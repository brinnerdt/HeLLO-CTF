module low_1 ( inData, clk, reset, outData );
  input [31:0] inData;
  output [31:0] outData;
  input clk, reset;
  wire   n23829, n23686, n23840, n23885, n12452, _________________18785,
         _________9_______18814, n23668, n23898, n12587, n12558, n12517,
         n23878, n23877, n23773, n23786, n12487, n23861, n23869, n23864,
         n12473, n12376, ______9__34498, n12413, n23946, n23945, n12511,
         n12346, n23941, n23942, n23943, n23909, __________0_____, n12520,
         n23669, n12478, n12442, n23920, __________0_______18820, n23704,
         _____9___34413, n23936, ______0__34499, n12412, n23801, n23882,
         n23924, n12547, _____9___34419, n23706, n12440, n23851, n23799,
         n23803, n23884, n23937, _____90__34411, __________0_______18822,
         n23772, n23800, n12522, n23997, n12564, n12384, n24032, n24024,
         n24026, n24035, n24030, n24025, n24023, n24028, n24027, n24029,
         n24033, n24031, n23850, n23922, n23672, n12414, n23928, n23671,
         n12402, n12310, n12371, n23903, n23991, n23831, n23845, n23782,
         n23788, n23789, n23856, n23859, n23814, n23715, n23857, n23767,
         n23865, n23867, n23969, n12297, n23960, n23971, n12506, n12330,
         n23712, n23860, n24045, n12546, n12515, n23921, n12580,
         __________0_______18819, n12391, n23667, __________0_______18818,
         n12426, n23681, n23797, n23804, n12476, n23995, n24021, n23979,
         n24012, n24002, n24003, n23982, n24020, n24013, n23983, n23972,
         n23992, n24001, n24008, n23990, n23999, n23998, n23970, n24009,
         n24000, n23964, n24006, n23963, n23974, n24007, n23962, n23976,
         n24004, n23975, n23978, n23977, n24005, n24038, n24039, n12316,
         n12472, n12355, n24042, n24046, n24040, n24047, n23986, n24017,
         n24055, n24051, n23871, n23872, n23837, n23893, n24037, n23873,
         n23894, n23895, n23836, n23892, n24036, n23838, n24057, n24048,
         n24062, n24053, n24059, n24052, n24061, n24056, n24054, n24058,
         n12464, n12408, n12331, n24019, n24015, n12393, n12340, n23958,
         n12333, n23993, n24011, n24022, n23948, n12302, n12319, n23959,
         n12299, n12320, n23951, n23953, n12388, n12305, n12401, n12586,
         n23985, n23981, n12394, n23828, n23987, n12392, n23949, n23950,
         n23938, n12380, n23961, n12584, n23932, n12373, n23705, n12484,
         n12429, n12513, n23740, n23760, n23741, n23728, n23727, n12479,
         n23693, n23763, n23738, n23694, n23762, n23720, n23737, n23765,
         n23736, n23875, n23876, n23833, n12450, n23843, n23711, n12451,
         n12486, n12583, n12481, n23754, n23725, n23682, n12480, n23745,
         n23753, n12475, n23757, n23746, n23747, n23748, n12441, n23756,
         n23683, n23733, n23742, n23743, n23758, n23730, n12516, n23830,
         n12430, n23848, n23853, n23714, n23854, n12518, n23880, n23750,
         n12351, n23759, n12485, n23793, n23697, n12446, n12445, n12521,
         n12549, n12354, n23666, n23774, n23775, n23783, n23778, n23784,
         n23779, n12579, n23795, n23787, n23766, n23796, n23781, n23696,
         n23691, n23780, n12544, n23794, n23679, n23791, n23790,
         __________0___0___18817, n12308, n23858, n12482, n23808, n23809,
         n23811, n12581, n23826, n12582, n23676, n23702, n12510, n23687,
         n23709, n23863, n12372, n23815, n23925, n23770, n23680, n23721,
         n23769, n23870, n12467, n23934, n23935, n12318, n1, n2, n3, n4, n5,
         n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20,
         n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62,
         n63, n64, n65, n66, n67, n68, n69, n70, n198, n209, n215, n698, n755,
         n756, n769, n771, n779, n811, n818, n821, n1144, n1519, n1520, n1678,
         n1965, n2029, n2045, n2046, n2047, n2056, n2074, n2113, n2116, n2122,
         n10140, n10141, n10142, n10143, n10144, n10145, n10146, n10147,
         n10148, n10149, n10150, n10151, n10152, n10153, n10154, n10155,
         n10156, n10157, n10158, n10159, n10160, n10161, n10162, n10163,
         n10164, n10165, n10166, n10167, n10168, n10169, n10170, n10171,
         n10172, n10173, n10174, n10175, n10176, n10177, n10178, n10179,
         n10180, n10181, n10182, n10183, n10184, n10185, n10186, n10187,
         n10188, n10189, n10190, n10191, n10192, n10193, n10194, n10195,
         n10196, n10197, n10198, n10199, n10200, n10201, n10202, n10203,
         n10204, n10205, n10206, n10207, n10208, n10209, n10210, n10211,
         n10212, n10213, n10214, n10215, n10216, n10217, n10218, n10219,
         n10220, n10221, n10222, n10223, n10224, n10225, n10226, n10227,
         n10228, n10229, n10230, n10231, n10232, n10233, n10234, n10235,
         n10236, n10237, n10238, n10239, n10240, n10241, n10242, n10243,
         n10244, n10245, n10246, n10247, n10248, n10249, n10250, n10251,
         n10252, n10253, n10254, n10255, n10256, n10257, n10258, n10259,
         n10260, n10261, n10262, n10263, n10264, n10265, n10266, n10267,
         n10268, n10269, n10270, n10271, n10272, n10273, n10274, n10275,
         n10276, n10277, n10278, n10279, n10280, n10281, n10282, n10283,
         n10284, n10285, n10286, n10287, n10288, n10289, n10290, n10291,
         n10292, n10293, n10294, n10295, n10296, n10297, n10298, n10299,
         n10300, n10301, n10302, n10303, n10304, n10305, n10306, n10307,
         n10308, n10309, n10310, n10311, n10312, n10313, n10314, n10315,
         n10316, n10317, n10318, n10319, n10320, n10321, n10322, n10323,
         n10324, n10325, n10326, n10327, n10328, n10329, n10330, n10331,
         n10332, n10333, n10334, n10335, n10336, n10337, n10338, n10339,
         n10340, n10341, n10342, n10343, n10344, n10345, n10346, n10347,
         n10348, n10349, n10350, n10351, n10352, n10353, n10354, n10355,
         n10356, n10357, n10358, n10359, n10360, n10361, n10362, n10363,
         n10364, n10365, n10366, n10367, n10368, n10369, n10370, n10371,
         n10372, n10373, n10374, n10375, n10376, n10377, n10378, n10379,
         n10380, n10381, n10382, n10383, n10384, n10385, n10386, n10387,
         n10388, n10389, n10390, n10391, n10392, n10393, n10394, n10395,
         n10396, n10397, n10398, n10399, n10400, n10401, n10402, n10403,
         n10404, n10405, n10406, n10407, n10408, n10409, n10410, n10411,
         n10412, n10413, n10414, n10415, n10416, n10417, n10418, n10419,
         n10420, n10421, n10422, n10423, n10424, n10425, n10426, n10427,
         n10428, n10429, n10430, n10431, n10432, n10433, n10434, n10435,
         n10436, n10437, n10438, n10439, n10440, n10441, n10442, n10443,
         n10444, n10445, n10446, n10447, n10448, n10449, n10450, n10451,
         n10452, n10453, n10454, n10455, n10456, n10457, n10458, n10459,
         n10460, n10461, n10462, n10463, n10464, n10465, n10466, n10467,
         n10468, n10469, n10470, n10471, n10472, n10473, n10474, n10475,
         n10476, n10477, n10478, n10479, n10480, n10481, n10482, n10483,
         n10484, n10485, n10486, n10487, n10488, n10489, n10490, n10491,
         n10492, n10493, n10494, n10495, n10496, n10497, n10498, n10499,
         n10500, n10501, n10502, n10503, n10504, n10505, n10506, n10507,
         n10508, n10509, n10510, n10511, n10512, n10513, n10514, n10515,
         n10516, n10517, n10518, n10519, n10520, n10521, n10522, n10523,
         n10524, n10525, n10526, n10527, n10528, n10529, n10530, n10531,
         n10532, n10533, n10534, n10535, n10536, n10537, n10538, n10539,
         n10540, n10541, n10542, n10543, n10544, n10545, n10546, n10547,
         n10548, n10549, n10550, n10551, n10552, n10553, n10554, n10555,
         n10556, n10557, n10558, n10559, n10560, n10561, n10562, n10563,
         n10564, n10565, n10566, n10567, n10568, n10569, n10570, n10571,
         n10572, n10573, n10574, n10575, n10576, n10577, n10578, n10579,
         n10580, n10581, n10582, n10583, n10584, n10585, n10586, n10587,
         n10588, n10589, n10590, n10591, n10592, n10593, n10594, n10595,
         n10596, n10597, n10598, n10599, n10600, n10601, n10602, n10603,
         n10604, n10605, n10606, n10607, n10608, n10609, n10610, n10611,
         n10612, n10613, n10614, n10615, n10616, n10617, n10618, n10619,
         n10620, n10621, n10622, n10623, n10624, n10625, n10626, n10627,
         n10628, n10629, n10630, n10631, n10632, n10633, n10634, n10635,
         n10636, n10637, n10638, n10639, n10640, n10641, n10642, n10643,
         n10644, n10645, n10646, n10647, n10648, n10649, n10650, n10651,
         n10652, n10653, n10654, n10655, n10656, n10657, n10658, n10659,
         n10660, n10661, n10662, n10663, n10664, n10665, n10666, n10667,
         n10668, n10669, n10670, n10671, n10672, n10673, n10674, n10675,
         n10676, n10677, n10678, n10679, n10680, n10681, n10682, n10683,
         n10684, n10685, n10686, n10687, n10688, n10689, n10690, n10691,
         n10692, n10693, n10694, n10695, n10696, n10697, n10698, n10699,
         n10700, n10701, n10702, n10703, n10704, n10705, n10706, n10707,
         n10708, n10709, n10710, n10711, n10712, n10713, n10714, n10715,
         n10716, n10717, n10718, n10719, n10720, n10721, n10722, n10723,
         n10724, n10725, n10726, n10727, n10728, n10729, n10730, n10731,
         n10732, n10733, n10734, n10735, n10736, n10737, n10738, n10739,
         n10740, n10741, n10742, n10743, n10744, n10745, n10746, n10747,
         n10748, n10749, n10750, n10751, n10752, n10753, n10754, n10755,
         n10756, n10757, n10758, n10759, n10760, n10761, n10762, n10763,
         n10764, n10765, n10766, n10767, n10768, n10769, n10770, n10771,
         n10772, n10773, n10774, n10775, n10776, n10777, n10778, n10779,
         n10780, n10781, n10782, n10783, n10784, n10785, n10786, n10787,
         n10788, n10789, n10790, n10791, n10792, n10793, n10794, n10795,
         n10796, n10797, n10798, n10799, n10800, n10801, n10802, n10803,
         n10804, n10805, n10806, n10807, n10808, n10809, n10810, n10811,
         n10812, n10813, n10814, n10815, n10816, n10817, n10818, n10819,
         n10820, n10821, n10822, n10823, n10824, n10825, n10826, n10827,
         n10828, n10829, n10830, n10831, n10832, n10833, n10834, n10835,
         n10836, n10837, n10838, n10839, n10840, n10841, n10842, n10843,
         n10844, n10845, n10846, n10847, n10848, n10849, n10850, n10851,
         n10852, n10853, n10854, n10855, n10856, n10857, n10858, n10859,
         n10860, n10861, n10862, n10863, n10864, n10865, n10866, n10867,
         n10868, n10869, n10870, n10871, n10872, n10873, n10874, n10875,
         n10876, n10877, n10878, n10879, n10880, n10881, n10882, n10883,
         n10884, n10885, n10886, n10887, n10888, n10889, n10890, n10891,
         n10892, n10893, n10894, n10895, n10896, n10897, n10898, n10899,
         n10900, n10901, n10902, n10903, n10904, n10905, n10906, n10907,
         n10908, n10909, n10910, n10911, n10912, n10913, n10914, n10915,
         n10916, n10917, n10918, n10919, n10920, n10921, n10922, n10923,
         n10924, n10925, n10926, n10927, n10928, n10929, n10930, n10931,
         n10932, n10933, n10934, n10935, n10936, n10937, n10938, n10939,
         n10940, n10941, n10942, n10943, n10944, n10945, n10946, n10947,
         n10948, n10949, n10950, n10951, n10952, n10953, n10954, n10955,
         n10956, n10957, n10958, n10959, n10960, n10961, n10962, n10963,
         n10964, n10965, n10966, n10967, n10968, n10969, n10970, n10971,
         n10972, n10973, n10974, n10975, n10976, n10977, n10978, n10979,
         n10980, n10981, n10982, n10983, n10984, n10985, n10986, n10987,
         n10988, n10989, n10990, n10991, n10992, n10993, n10994, n10995,
         n10996, n10997, n10998, n10999, n11000, n11001, n11002, n11003,
         n11004, n11005, n11006, n11007, n11008, n11009, n11010, n11011,
         n11012, n11013, n11014, n11015, n11016, n11017, n11018, n11019,
         n11020, n11021, n11022, n11023, n11024, n11025, n11026, n11027,
         n11028, n11029, n11030, n11031, n11032, n11033, n11034, n11035,
         n11036, n11037, n11038, n11039, n11040, n11041, n11042, n11043,
         n11044, n11045, n11046, n11047, n11048, n11049, n11050, n11051,
         n11052, n11053, n11054, n11055, n11056, n11057, n11058, n11059,
         n11060, n11061, n11062, n11063, n11064, n11065, n11066, n11067,
         n11068, n11069, n11070, n11071, n11072, n11073, n11074, n11075,
         n11076, n11077, n11078, n11079, n11080, n11081, n11082, n11083,
         n11084, n11085, n11086, n11087, n11088, n11089, n11090, n11091,
         n11092, n11093, n11094, n11095, n11096, n11097, n11098, n11099,
         n11100, n11101, n11102, n11103, n11104, n11105, n11106, n11107,
         n11108, n11109, n11110, n11111, n11112, n11113, n11114, n11115,
         n11116, n11117, n11118, n11119, n11120, n11121, n11122, n11123,
         n11124, n11125, n11126, n11127, n11128, n11129, n11130, n11131,
         n11132, n11133, n11134, n11135, n11136, n11137, n11138, n11139,
         n11140, n11141, n11142, n11143, n11144, n11145, n11146, n11147,
         n11148, n11149, n11150, n11151, n11152, n11153, n11154, n11155,
         n11156, n11157, n11158, n11159, n11160, n11161, n11162, n11163,
         n11164, n11165, n11166, n11167, n11168, n11169, n11170, n11171,
         n11172, n11173, n11174, n11175, n11176, n11177, n11178, n11179,
         n11180, n11181, n11182, n11183, n11184, n11185, n11186, n11187,
         n11188, n11189, n11190, n11191, n11192, n11193, n11194, n11195,
         n11196, n11197, n11198, n11199, n11200, n11201, n11202, n11203,
         n11204, n11205, n11206, n11207, n11208, n11209, n11210, n11211,
         n11212, n11213, n11214, n11215, n11216, n11217, n11218, n11219,
         n11220, n11221, n11222, n11223, n11224, n11225, n11226, n11227,
         n11228, n11229, n11230, n11231, n11232, n11233, n11234, n11235,
         n11236, n11237, n11238, n11239, n11240, n11241, n11242, n11243,
         n11244, n11245, n11246, n11247, n11248, n11249, n11250, n11251,
         n11252, n11253, n11254, n11255, n11256, n11257, n11258, n11259,
         n11260, n11261, n11262, n11263, n11264, n11265, n11266, n11267,
         n11268, n11269, n11270, n11271, n11272, n11273, n11274, n11275,
         n11276, n11277, n11278, n11279, n11280, n11281, n11282, n11283,
         n11284, n11285, n11286, n11287, n11288, n11289, n11290, n11291,
         n11292, n11293, n11294, n11295, n11296, n11297, n11298, n11299,
         n11300, n11301, n11302, n11303, n11304, n11305, n11306, n11307,
         n11308, n11309, n11310, n11311, n11312, n11313, n11314, n11315,
         n11316, n11317, n11318, n11319, n11320, n11321, n11322, n11323,
         n11324, n11325, n11326, n11327, n11328, n11329, n11330, n11331,
         n11332, n11333, n11334, n11335, n11336, n11337, n11338, n11339,
         n11340, n11341, n11342, n11343, n11344, n11345, n11346, n11347,
         n11348, n11349, n11350, n11351, n11352, n11353, n11354, n11355,
         n11356, n11357, n11358, n11359, n11360, n11361, n11362, n11363,
         n11364, n11365, n11366, n11367, n11368, n11369, n11370, n11371,
         n11372, n11373, n11374, n11375, n11376, n11377, n11378, n11379,
         n11380, n11381, n11382, n11383, n11384, n11385, n11386, n11387,
         n11388, n11389, n11390, n11391, n11392, n11393, n11394, n11395,
         n11396, n11397, n11398, n11399, n11400, n11401, n11402, n11403,
         n11404, n11405, n11406, n11407, n11408, n11409, n11410, n11411,
         n11412, n11413, n11414, n11415, n11416, n11417, n11418, n11419,
         n11420, n11421, n11422, n11423, n11424, n11425, n11426, n11427,
         n11428, n11429, n11430, n11431, n11432, n11433, n11434, n11435,
         n11436, n11437, n11438, n11439, n11440, n11441, n11442, n11443,
         n11444, n11445, n11446, n11447, n11448, n11449, n11450, n11451,
         n11452, n11453, n11454, n11455, n11456, n11457, n11458, n11459,
         n11460, n11461, n11462, n11463, n11464, n11465, n11466, n11467,
         n11468, n11469, n11470, n11471, n11472, n11473, n11474, n11475,
         n11476, n11477, n11478, n11479, n11480, n11481, n11482, n11483,
         n11484, n11485, n11486, n11487, n11488, n11489, n11490, n11491,
         n11492, n11493, n11494, n11495, n11496, n11497, n11498, n11499,
         n11500, n11501, n11502, n11503, n11504, n11505, n11506, n11507,
         n11508, n11509, n11510, n11511, n11512, n11513, n11514, n11515,
         n11516, n11517, n11518, n11519, n11520, n11521, n11522, n11523,
         n11524, n11525, n11526, n11527, n11528, n11529, n11530, n11531,
         n11532, n11533, n11534, n11535, n11536, n11537, n11538, n11539,
         n11540, n11541, n11542, n11543, n11544, n11545, n11546, n11547,
         n11548, n11549, n11550, n11551, n11552, n11553, n11554, n11555,
         n11556, n11557, n11558, n11559, n11560, n11561, n11562, n11563,
         n11564, n11565, n11566, n11567, n11568, n11569, n11570, n11571,
         n11572, n11573, n11574, n11575, n11576, n11577, n11578, n11579,
         n11580, n11581, n11582, n11583, n11584, n11585, n11586, n11587,
         n11588, n11589, n11590, n11591, n11592, n11593, n11594, n11595,
         n11596, n11597, n11598, n11599, n11600, n11601, n11602, n11603,
         n11604, n11605, n11606, n11607, n11608, n11609, n11610, n11611,
         n11612, n11613, n11614, n11615, n11616, n11617, n11618, n11619,
         n11620, n11621, n11622, n11623, n11624, n11625, n11626, n11627,
         n11628, n11629, n11630, n11631, n11632, n11633, n11634, n11635,
         n11636, n11637, n11638, n11639, n11640, n11641, n11642, n11643,
         n11644, n11645, n11646, n11647, n11648, n11649, n11650, n11651,
         n11652, n11653, n11654, n11655, n11656, n11657, n11658, n11659,
         n11660, n11661, n11662, n11663, n11664, n11665, n11666, n11667,
         n11668, n11669, n11670, n11671, n11672, n11673, n11674, n11675,
         n11676, n11677, n11678, n11679, n11680, n11681, n11682, n11683,
         n11684, n11685, n11686, n11687, n11688, n11689, n11690, n11691,
         n11692, n11693, n11694, n11695, n11696, n11697, n11698, n11699,
         n11700, n11701, n11702, n11703, n11704, n11705, n11706, n11707,
         n11708, n11709, n11710, n11711, n11712, n11713, n11714, n11715,
         n11716, n11717, n11718, n11719, n11720, n11721, n11722, n11723,
         n11724, n11725, n11726, n11727, n11728, n11729, n11730, n11731,
         n11732, n11733, n11734, n11735, n11736, n11737, n11738, n11739,
         n11740, n11741, n11742, n11743, n11744, n11745, n11746, n11747,
         n11748, n11749, n11750, n11751, n11752, n11753, n11754, n11755,
         n11756, n11757, n11758, n11759, n11760, n11761, n11762, n11763,
         n11764, n11765, n11766, n11767, n11768, n11769, n11770, n11771,
         n11772, n11773, n11774, n11775, n11776, n11777, n11778, n11779,
         n11780, n11781, n11782, n11783, n11784, n11785, n11786, n11787,
         n11788, n11789, n11790, n11791, n11792, n11793, n11794, n11795,
         n11796, n11797, n11798, n11799, n11800, n11801, n11802, n11803,
         n11804, n11805, n11806, n11807, n11808, n11809, n11810, n11811,
         n11812, n11813, n11814, n11815, n11816, n11817, n11818, n11819,
         n11820, n11821, n11822, n11823, n11824, n11825, n11826, n11827,
         n11828, n11829, n11830, n11831, n11832, n11833, n11834, n11835,
         n11836, n11837, n11838, n11839, n11840, n11841, n11842, n11843,
         n11844, n11845, n11846, n11847, n11848, n11849, n11850, n11851,
         n11852, n11853, n11854, n11855, n11856, n11857, n11858, n11859,
         n11860, n11861, n11862, n11863, n11864, n11865, n11866, n11867,
         n11868, n11869, n11870, n11871, n11872, n11873, n11874, n11875,
         n11876, n11877, n11878, n11879, n11880, n11881, n11882, n11883,
         n11884, n11885, n11886, n11887, n11888, n11889, n11890, n11891,
         n11892, n11893, n11894, n11895, n11896, n11897, n11898, n11899,
         n11900, n11901, n11902, n11903, n11904, n11905, n11906, n11907,
         n11908, n11909, n11910, n11911, n11912, n11913, n11914, n11915,
         n11916, n11917, n11918, n11919, n11920, n11921, n11922, n11923,
         n11924, n11925, n11926, n11927, n11928, n11929, n11930, n11931,
         n11932, n11933, n11934, n11935, n11936, n11937, n11938, n11939,
         n11940, n11941, n11942, n11943, n11944, n11945, n11946, n11947,
         n11948, n11949, n11950, n11951, n11952, n11953, n11954, n11955,
         n11956, n11957, n11958, n11959, n11960, n11961, n11962, n11963,
         n11964, n11965, n11966, n11967, n11968, n11969, n11970, n11971,
         n11972, n11973, n11974, n11975, n11976, n11977, n11978, n11979,
         n11980, n11981, n11982, n11983, n11984, n11985, n11986, n11987,
         n11988, n11989, n11990, n11991, n11992, n11993, n11994, n11995,
         n11996, n11997, n11998, n11999, n12000, n12001, n12002, n12003,
         n12004, n12005, n12006, n12007, n12008, n12009, n12010, n12011,
         n12012, n12013, n12014, n12015, n12016, n12017, n12018, n12019,
         n12020, n12021, n12022, n12023, n12024, n12025, n12026, n12027,
         n12028, n12029, n12030, n12031, n12032, n12033, n12034, n12035,
         n12036, n12037, n12038, n12039, n12040, n12041, n12042, n12043,
         n12044, n12045, n12046, n12047, n12048, n12049, n12050, n12051,
         n12052, n12053, n12054, n12055, n12056, n12057, n12058, n12059,
         n12060, n12061, n12062, n12063, n12064, n12065, n12066, n12067,
         n12068, n12069, n12070, n12071, n12072, n12073, n12074, n12075,
         n12076, n12077, n12078, n12079, n12080, n12081, n12082, n12083,
         n12084, n12085, n12086, n12087, n12088, n12089, n12090, n12091,
         n12092, n12093, n12094, n12095, n12096, n12097, n12098, n12099,
         n12100, n12101, n12102, n12103, n12104, n12105, n12106, n12107,
         n12108, n12109, n12110, n12111, n12112, n12113, n12114, n12115,
         n12116, n12117, n12118, n12119, n12120, n12121, n12122, n12123,
         n12124, n12125, n12126, n12127, n12128, n12129, n12130, n12131,
         n12132, n12133, n12134, n12135, n12136, n12137, n12138, n12139,
         n12140, n12141, n12142, n12143, n12144, n12145, n12146, n12147,
         n12148, n12149, n12150, n12151, n12152, n12153, n12154, n12155,
         n12156, n12157, n12158, n12159, n12160, n12161, n12162, n12163,
         n12164, n12165, n12166, n12167, n12168, n12169, n12170, n12171,
         n12172, n12173, n12174, n12175, n12176, n12177, n12178, n12179,
         n12180, n12181, n12182, n12183, n12184, n12185, n12186, n12187,
         n12188, n12189, n12190, n12191, n12192, n12193, n12194, n12195,
         n12196, n12197, n12198, n12199, n12200, n12201, n12202, n12203,
         n12204, n12205, n12206, n12207, n12208, n12209, n12210, n12211,
         n12212, n12213, n12214, n12215, n12216, n12217, n12218, n12219,
         n12220, n12221, n12222, n12223, n12224, n12225, n12226, n12227,
         n12228, n12229, n12230, n12231, n12232, n12233, n12234, n12235,
         n12236, n12237, n12238, n12239, n12240, n12241, n12242, n12243,
         n12244, n12245, n12246, n12247, n12248, n12249, n12250, n12251,
         n12252, n12253, n12254, n12255, n12256, n12257, n12258, n12259,
         n12260, n12261, n12262, n12263, n12264, n12265, n12266, n12267,
         n12268, n12269, n12270, n12271, n12272, n12273, n12274, n12275,
         n12276, n12277, n12278, n12279, n12280, n12281, n12282, n12283,
         n12284, n12285, n12286, n12287, n12288, n12289, n12290, n12291,
         n12292, n12293, n12294, n12295, n12296, n12298, n12300, n12301,
         n12303, n12304, n12306, n12307, n12309, n12311, n12312, n12313,
         n12314, n12315, n12317, n12321, n12322, n12323, n12324, n12325,
         n12326, n12327, n12328, n12329, n12332, n12334, n12335, n12336,
         n12337, n12338, n12339, n12341, n12342, n12343, n12344, n12345,
         n12347, n12348, n12349, n12350, n12352, n12353, n12356, n12357,
         n12358, n12359, n12360, n12361, n12362, n12363, n12364, n12365,
         n12366, n12367, n12368, n12369, n12370, n12374, n12375, n12377,
         n12378, n12379, n12381, n12382, n12383, n12385, n12386, n12387,
         n12389, n12390, n12395, n12396, n12397, n12398, n12399, n12400,
         n12403, n12404, n12405, n12406, n12407, n12409, n12410, n12411,
         n12415, n12416, n12417, n12418, n12419, n12420, n12421, n12422,
         n12423, n12424, n12425, n12427, n12428, n12431, n12432, n12433,
         n12434, n12435, n12436, n12437, n12438, n12439, n12443, n12444,
         n12447, n12448, n12449, n12453, n12454, n12455, n12456, n12457,
         n12458, n12459, n12460, n12461, n12462, n12463, n12465, n12466,
         n12468, n12469, n12470, n12471, n12474, n12477, n12483, n12488,
         n12489, n12490, n12491, n12492, n12493, n12494, n12495, n12496,
         n12497, n12498, n12499, n12500, n12501, n12502, n12503, n12504,
         n12505, n12507, n12508, n12509, n12512, n12514, n12519, n12523,
         n12524, n12525, n12526, n12527, n12528, n12529, n12530, n12531,
         n12532, n12533, n12534, n12535, n12536, n12537, n12538, n12539,
         n12540, n12541, n12542, n12543, n12545, n12548, n12550, n12551,
         n12552, n12553, n12554, n12555, n12556, n12557, n12559, n12560,
         n12561, n12562, n12563, n12565, n12566, n12567, n12568, n12569,
         n12570, n12571, n12572, n12573, n12574, n12575, n12576, n12577,
         n12578, n12585, n12588, n12589, n12590, n12591, n12592, n12593,
         n12594, n12595, n12596, n12597, n12598, n12599, n12600, n12601,
         n12602, n12603, n12604, n12605, n12606, n12607, n12608, n12609,
         n12610, n12611, n12612, n12613, n12614, n12615, n12616, n12617,
         n12618, n12619, n12620, n12621, n12622, n12623, n12624, n12625,
         n12626, n12627, n12628, n12629, n12630, n12631, n12632, n12633,
         n12634, n12635, n12636, n12637, n12638, n12639, n12640, n12641,
         n12642, n12643, n12644, n12645, n12646, n12647, n12648, n12649,
         n12650, n12651, n12652, n12653, n12654, n12655, n12656, n12657,
         n12658, n12659, n12660, n12661, n12662, n12663, n12664, n12665,
         n12666, n12667, n12668, n12669, n12670, n12671, n12672, n12673,
         n12674, n12675, n12676, n12677, n12678, n12679, n12680, n12681,
         n12682, n12683, n12684, n12685, n12686, n12687, n12688, n12689,
         n12690, n12691, n12692, n12693, n12694, n12695, n12696, n12697,
         n12698, n12699, n12700, n12701, n12702, n12703, n12704, n12705,
         n12706, n12707, n12708, n12709, n12710, n12711, n12712, n12713,
         n12714, n12715, n12716, n12717, n12718, n12719, n12720, n12721,
         n12722, n12723, n12724, n12725, n12726, n12727, n12728, n12729,
         n12730, n12731, n12732, n12733, n12734, n12735, n12736, n12737,
         n12738, n12739, n12740, n12741, n12742, n12743, n12744, n12745,
         n12746, n12747, n12748, n12749, n12750, n12751, n12752, n12753,
         n12754, n12755, n12756, n12757, n12758, n12759, n12760, n12761,
         n12762, n12763, n12764, n12765, n12766, n12767, n12768, n12769,
         n12770, n12771, n12772, n12773, n12774, n12775, n12776, n12777,
         n12778, n12779, n12780, n12781, n12782, n12783, n12784, n12785,
         n12786, n12787, n12788, n12789, n12790, n12791, n12792, n12793,
         n12794, n12795, n12796, n12797, n12798, n12799, n12800, n12801,
         n12802, n12803, n12804, n12805, n12806, n12807, n12808, n12809,
         n12810, n12811, n12812, n12813, n12814, n12815, n12816, n12817,
         n12818, n12819, n12820, n12821, n12822, n12823, n12824, n12825,
         n12826, n12827, n12828, n12829, n12830, n12831, n12832, n12833,
         n12834, n12835, n12836, n12837, n12838, n12839, n12840, n12841,
         n12842, n12843, n12844, n12845, n12846, n12847, n12848, n12849,
         n12850, n12851, n12852, n12853, n12854, n12855, n12856, n12857,
         n12858, n12859, n12860, n12861, n12862, n12863, n12864, n12865,
         n12866, n12867, n12868, n12869, n12870, n12871, n12872, n12873,
         n12874, n12875, n12876, n12877, n12878, n12879, n12880, n12881,
         n12882, n12883, n12884, n12885, n12886, n12887, n12888, n12889,
         n12890, n12891, n12892, n12893, n12894, n12895, n12896, n12897,
         n12898, n12899, n12900, n12901, n12902, n12903, n12904, n12905,
         n12906, n12907, n12908, n12909, n12910, n12911, n12912, n12913,
         n12914, n12915, n12916, n12917, n12918, n12919, n12920, n12921,
         n12922, n12923, n12924, n12925, n12926, n12927, n12928, n12929,
         n12930, n12931, n12932, n12933, n12934, n12935, n12936, n12937,
         n12938, n12939, n12940, n12941, n12942, n12943, n12944, n12945,
         n12946, n12947, n12948, n12949, n12950, n12951, n12952, n12953,
         n12954, n12955, n12956, n12957, n12958, n12959, n12960, n12961,
         n12962, n12963, n12964, n12965, n12966, n12967, n12968, n12969,
         n12970, n12971, n12972, n12973, n12974, n12975, n12976, n12977,
         n12978, n12979, n12980, n12981, n12982, n12983, n12984, n12985,
         n12986, n12987, n12988, n12989, n12990, n12991, n12992, n12993,
         n12994, n12995, n12996, n12997, n12998, n12999, n13000, n13001,
         n13002, n13003, n13004, n13005, n13006, n13007, n13008, n13009,
         n13010, n13011, n13012, n13013, n13014, n13015, n13016, n13017,
         n13018, n13019, n13020, n13021, n13022, n13023, n13024, n13025,
         n13026, n13027, n13028, n13029, n13030, n13031, n13032, n13033,
         n13034, n13035, n13036, n13037, n13038, n13039, n13040, n13041,
         n13042, n13043, n13044, n13045, n13046, n13047, n13048, n13049,
         n13050, n13051, n13052, n13053, n13054, n13055, n13056, n13057,
         n13058, n13059, n13060, n13061, n13062, n13063, n13064, n13065,
         n13066, n13067, n13068, n13069, n13070, n13071, n13072, n13073,
         n13074, n13075, n13076, n13077, n13078, n13079, n13080, n13081,
         n13082, n13083, n13084, n13085, n13086, n13087, n13088, n13089,
         n13090, n13091, n13092, n13093, n13094, n13095, n13096, n13097,
         n13098, n13099, n13100, n13101, n13102, n13103, n13104, n13105,
         n13106, n13107, n13108, n13109, n13110, n13111, n13112, n13113,
         n13114, n13115, n13116, n13117, n13118, n13119, n13120, n13121,
         n13122, n13123, n13124, n13125, n13126, n13127, n13128, n13129,
         n13130, n13131, n13132, n13133, n13134, n13135, n13136, n13137,
         n13138, n13139, n13140, n13141, n13142, n13143, n13144, n13145,
         n13146, n13147, n13148, n13149, n13150, n13151, n13152, n13153,
         n13154, n13155, n13156, n13157, n13158, n13159, n13160, n13161,
         n13162, n13163, n13164, n13165, n13166, n13167, n13168, n13169,
         n13170, n13171, n13172, n13173, n13174, n13175, n13176, n13177,
         n13178, n13179, n13180, n13181, n13182, n13183, n13184, n13185,
         n13186, n13187, n13188, n13189, n13190, n13191, n13192, n13193,
         n13194, n13195, n13196, n13197, n13198, n13199, n13200, n13201,
         n13202, n13203, n13204, n13205, n13206, n13207, n13208, n13209,
         n13210, n13211, n13212, n13213, n13214, n13215, n13216, n13217,
         n13218, n13219, n13220, n13221, n13222, n13223, n13224, n13225,
         n13226, n13227, n13228, n13229, n13230, n13231, n13232, n13233,
         n13234, n13235, n13236, n13237, n13238, n13239, n13240, n13241,
         n13242, n13243, n13244, n13245, n13246, n13247, n13248, n13249,
         n13250, n13251, n13252, n13253, n13254, n13255, n13256, n13257,
         n13258, n13259, n13260, n13261, n13262, n13263, n13264, n13265,
         n13266, n13267, n13268, n13269, n13270, n13271, n13272, n13273,
         n13274, n13275, n13276, n13277, n13278, n13279, n13280, n13281,
         n13282, n13283, n13284, n13285, n13286, n13287, n13288, n13289,
         n13290, n13291, n13292, n13293, n13294, n13295, n13296, n13297,
         n13298, n13299, n13300, n13301, n13302, n13303, n13304, n13305,
         n13306, n13307, n13308, n13309, n13310, n13311, n13312, n13313,
         n13314, n13315, n13316, n13317, n13318, n13319, n13320, n13321,
         n13322, n13323, n13324, n13325, n13326, n13327, n13328, n13329,
         n13330, n13331, n13332, n13333, n13334, n13335, n13336, n13337,
         n13338, n13339, n13340, n13341, n13342, n13343, n13344, n13345,
         n13346, n13347, n13348, n13349, n13350, n13351, n13352, n13353,
         n13354, n13355, n13356, n13357, n13358, n13359, n13360, n13361,
         n13362, n13363, n13364, n13365, n13366, n13367, n13368, n13369,
         n13370, n13371, n13372, n13373, n13374, n13375, n13376, n13377,
         n13378, n13379, n13380, n13381, n13382, n13383, n13384, n13385,
         n13386, n13387, n13388, n13389, n13390, n13391, n13392, n13393,
         n13394, n13395, n13396, n13397, n13398, n13399, n13400, n13401,
         n13402, n13403, n13404, n13405, n13406, n13407, n13408, n13409,
         n13410, n13411, n13412, n13413, n13414, n13415, n13416, n13417,
         n13418, n13419, n13420, n13421, n13422, n13423, n13424, n13425,
         n13426, n13427, n13428, n13429, n13430, n13431, n13432, n13433,
         n13434, n13435, n13436, n13437, n13438, n13439, n13440, n13441,
         n13442, n13443, n13444, n13445, n13446, n13447, n13448, n13449,
         n13450, n13451, n13452, n13453, n13454, n13455, n13456, n13457,
         n13458, n13459, n13460, n13461, n13462, n13463, n13464, n13465,
         n13466, n13467, n13468, n13469, n13470, n13471, n13472, n13473,
         n13474, n13475, n13476, n13477, n13478, n13479, n13480, n13481,
         n13482, n13483, n13484, n13485, n13486, n13487, n13488, n13489,
         n13490, n13491, n13492, n13493, n13494, n13495, n13496, n13497,
         n13498, n13499, n13500, n13501, n13502, n13503, n13504, n13505,
         n13506, n13507, n13508, n13509, n13510, n13511, n13512, n13513,
         n13514, n13515, n13516, n13517, n13518, n13519, n13520, n13521,
         n13522, n13523, n13524, n13525, n13526, n13527, n13528, n13529,
         n13530, n13531, n13532, n13533, n13534, n13535, n13536, n13537,
         n13538, n13539, n13540, n13541, n13542, n13543, n13544, n13545,
         n13546, n13547, n13548, n13549, n13550, n13551, n13552, n13553,
         n13554, n13555, n13556, n13557, n13558, n13559, n13560, n13561,
         n13562, n13563, n13564, n13565, n13566, n13567, n13568, n13569,
         n13570, n13571, n13572, n13573, n13574, n13575, n13576, n13577,
         n13578, n13579, n13580, n13581, n13582, n13583, n13584, n13585,
         n13586, n13587, n13588, n13589, n13590, n13591, n13592, n13593,
         n13594, n13595, n13596, n13597, n13598, n13599, n13600, n13601,
         n13602, n13603, n13604, n13605, n13606, n13607, n13608, n13609,
         n13610, n13611, n13612, n13613, n13614, n13615, n13616, n13617,
         n13618, n13619, n13620, n13621, n13622, n13623, n13624, n13625,
         n13626, n13627, n13628, n13629, n13630, n13631, n13632, n13633,
         n13634, n13635, n13636, n13637, n13638, n13639, n13640, n13641,
         n13642, n13643, n13644, n13645, n13646, n13647, n13648, n13649,
         n13650, n13651, n13652, n13653, n13654, n13655, n13656, n13657,
         n13658, n13659, n13660, n13661, n13662, n13663, n13664, n13665,
         n13666, n13667, n13668, n13669, n13670, n13671, n13672, n13673,
         n13674, n13675, n13676, n13677, n13678, n13679, n13680, n13681,
         n13682, n13683, n13684, n13685, n13686, n13687, n13688, n13689,
         n13690, n13691, n13692, n13693, n13694, n13695, n13696, n13697,
         n13698, n13699, n13700, n13701, n13702, n13703, n13704, n13705,
         n13706, n13707, n13708, n13709, n13710, n13711, n13712, n13713,
         n13714, n13715, n13716, n13717, n13718, n13719, n13720, n13721,
         n13722, n13723, n13724, n13725, n13726, n13727, n13728, n13729,
         n13730, n13731, n13732, n13733, n13734, n13735, n13736, n13737,
         n13738, n13739, n13740, n13741, n13742, n13743, n13744, n13745,
         n13746, n13747, n13748, n13749, n13750, n13751, n13752, n13753,
         n13754, n13755, n13756, n13757, n13758, n13759, n13760, n13761,
         n13762, n13763, n13764, n13765, n13766, n13767, n13768, n13769,
         n13770, n13771, n13772, n13773, n13774, n13775, n13776, n13777,
         n13778, n13779, n13780, n13781, n13782, n13783, n13784, n13785,
         n13786, n13787, n13788, n13789, n13790, n13791, n13792, n13793,
         n13794, n13795, n13796, n13797, n13798, n13799, n13800, n13801,
         n13802, n13803, n13804, n13805, n13806, n13807, n13808, n13809,
         n13810, n13811, n13812, n13813, n13814, n13815, n13816, n13817,
         n13818, n13819, n13820, n13821, n13822, n13823, n13824, n13825,
         n13826, n13827, n13828, n13829, n13830, n13831, n13832, n13833,
         n13834, n13835, n13836, n13837, n13838, n13839, n13840, n13841,
         n13842, n13843, n13844, n13845, n13846, n13847, n13848, n13849,
         n13850, n13851, n13852, n13853, n13854, n13855, n13856, n13857,
         n13858, n13859, n13860, n13861, n13862, n13863, n13864, n13865,
         n13866, n13867, n13868, n13869, n13870, n13871, n13872, n13873,
         n13874, n13875, n13876, n13877, n13878, n13879, n13880, n13881,
         n13882, n13883, n13884, n13885, n13886, n13887, n13888, n13889,
         n13890, n13891, n13892, n13893, n13894, n13895, n13896, n13897,
         n13898, n13899, n13900, n13901, n13902, n13903, n13904, n13905,
         n13906, n13907, n13908, n13909, n13910, n13911, n13912, n13913,
         n13914, n13915, n13916, n13917, n13918, n13919, n13920, n13921,
         n13922, n13923, n13924, n13925, n13926, n13927, n13928, n13929,
         n13930, n13931, n13932, n13933, n13934, n13935, n13936, n13937,
         n13938, n13939, n13940, n13941, n13942, n13943, n13944, n13945,
         n13946, n13947, n13948, n13949, n13950, n13951, n13952, n13953,
         n13954, n13955, n13956, n13957, n13958, n13959, n13960, n13961,
         n13962, n13963, n13964, n13965, n13966, n13967, n13968, n13969,
         n13970, n13971, n13972, n13973, n13974, n13975, n13976, n13977,
         n13978, n13979, n13980, n13981, n13982, n13983, n13984, n13985,
         n13986, n13987, n13988, n13989, n13990, n13991, n13992, n13993,
         n13994, n13995, n13996, n13997, n13998, n13999, n14000, n14001,
         n14002, n14003, n14004, n14005, n14006, n14007, n14008, n14009,
         n14010, n14011, n14012, n14013, n14014, n14015, n14016, n14017,
         n14018, n14019, n14020, n14021, n14022, n14023, n14024, n14025,
         n14026, n14027, n14028, n14029, n14030, n14031, n14032, n14033,
         n14034, n14035, n14036, n14037, n14038, n14039, n14040, n14041,
         n14042, n14043, n14044, n14045, n14046, n14047, n14048, n14049,
         n14050, n14051, n14052, n14053, n14054, n14055, n14056, n14057,
         n14058, n14059, n14060, n14061, n14062, n14063, n14064, n14065,
         n14066, n14067, n14068, n14069, n14070, n14071, n14072, n14073,
         n14074, n14075, n14076, n14077, n14078, n14079, n14080, n14081,
         n14082, n14083, n14084, n14085, n14086, n14087, n14088, n14089,
         n14090, n14091, n14092, n14093, n14094, n14095, n14096, n14097,
         n14098, n14099, n14100, n14101, n14102, n14103, n14104, n14105,
         n14106, n14107, n14108, n14109, n14110, n14111, n14112, n14113,
         n14114, n14115, n14116, n14117, n14118, n14119, n14120, n14121,
         n14122, n14123, n14124, n14125, n14126, n14127, n14128, n14129,
         n14130, n14131, n14132, n14133, n14134, n14135, n14136, n14137,
         n14138, n14139, n14140, n14141, n14142, n14143, n14144, n14145,
         n14146, n14147, n14148, n14149, n14150, n14151, n14152, n14153,
         n14154, n14155, n14156, n14157, n14158, n14159, n14160, n14161,
         n14162, n14163, n14164, n14165, n14166, n14167, n14168, n14169,
         n14170, n14171, n14172, n14173, n14174, n14175, n14176, n14177,
         n14178, n14179, n14180, n14181, n14182, n14183, n14184, n14185,
         n14186, n14187, n14188, n14189, n14190, n14191, n14192, n14193,
         n14194, n14195, n14196, n14197, n14198, n14199, n14200, n14201,
         n14202, n14203, n14204, n14205, n14206, n14207, n14208, n14209,
         n14210, n14211, n14212, n14213, n14214, n14215, n14216, n14217,
         n14218, n14219, n14220, n14221, n14222, n14223, n14224, n14225,
         n14226, n14227, n14228, n14229, n14230, n14231, n14232, n14233,
         n14234, n14235, n14236, n14237, n14238, n14239, n14240, n14241,
         n14242, n14243, n14244, n14245, n14246, n14247, n14248, n14249,
         n14250, n14251, n14252, n14253, n14254, n14255, n14256, n14257,
         n14258, n14259, n14260, n14261, n14262, n14263, n14264, n14265,
         n14266, n14267, n14268, n14269, n14270, n14271, n14272, n14273,
         n14274, n14275, n14276, n14277, n14278, n14279, n14280, n14281,
         n14282, n14283, n14284, n14285, n14286, n14287, n14288, n14289,
         n14290, n14291, n14292, n14293, n14294, n14295, n14296, n14297,
         n14298, n14299, n14300, n14301, n14302, n14303, n14304, n14305,
         n14306, n14307, n14308, n14309, n14310, n14311, n14312, n14313,
         n14314, n14315, n14316, n14317, n14318, n14319, n14320, n14321,
         n14322, n14323, n14324, n14325, n14326, n14327, n14328, n14329,
         n14330, n14331, n14332, n14333, n14334, n14335, n14336, n14337,
         n14338, n14339, n14340, n14341, n14342, n14343, n14344, n14345,
         n14346, n14347, n14348, n14349, n14350, n14351, n14352, n14353,
         n14354, n14355, n14356, n14357, n14358, n14359, n14360, n14361,
         n14362, n14363, n14364, n14365, n14366, n14367, n14368, n14369,
         n14370, n14371, n14372, n14373, n14374, n14375, n14376, n14377,
         n14378, n14379, n14380, n14381, n14382, n14383, n14384, n14385,
         n14386, n14387, n14388, n14389, n14390, n14391, n14392, n14393,
         n14394, n14395, n14396, n14397, n14398, n14399, n14400, n14401,
         n14402, n14403, n14404, n14405, n14406, n14407, n14408, n14409,
         n14410, n14411, n14412, n14413, n14414, n14415, n14416, n14417,
         n14418, n14419, n14420, n14421, n14422, n14423, n14424, n14425,
         n14426, n14427, n14428, n14429, n14430, n14431, n14432, n14433,
         n14434, n14435, n14436, n14437, n14438, n14439, n14440, n14441,
         n14442, n14443, n14444, n14445, n14446, n14447, n14448, n14449,
         n14450, n14451, n14452, n14453, n14454, n14455, n14456, n14457,
         n14458, n14459, n14460, n14461, n14462, n14463, n14464, n14465,
         n14466, n14467, n14468, n14469, n14470, n14471, n14472, n14473,
         n14474, n14475, n14476, n14477, n14478, n14479, n14480, n14481,
         n14482, n14483, n14484, n14485, n14486, n14487, n14488, n14489,
         n14490, n14491, n14492, n14493, n14494, n14495, n14496, n14497,
         n14498, n14499, n14500, n14501, n14502, n14503, n14504, n14505,
         n14506, n14507, n14508, n14509, n14510, n14511, n14512, n14513,
         n14514, n14515, n14516, n14517, n14518, n14519, n14520, n14521,
         n14522, n14523, n14524, n14525, n14526, n14527, n14528, n14529,
         n14530, n14531, n14532, n14533, n14534, n14535, n14536, n14537,
         n14538, n14539, n14540, n14541, n14542, n14543, n14544, n14545,
         n14546, n14547, n14548, n14549, n14550, n14551, n14552, n14553,
         n14554, n14555, n14556, n14557, n14558, n14559, n14560, n14561,
         n14562, n14563, n14564, n14565, n14566, n14567, n14568, n14569,
         n14570, n14571, n14572, n14573, n14574, n14575, n14576, n14577,
         n14578, n14579, n14580, n14581, n14582, n14583, n14584, n14585,
         n14586, n14587, n14588, n14589, n14590, n14591, n14592, n14593,
         n14594, n14595, n14596, n14597, n14598, n14599, n14600, n14601,
         n14602, n14603, n14604, n14605, n14606, n14607, n14608, n14609,
         n14610, n14611, n14612, n14613, n14614, n14615, n14616, n14617,
         n14618, n14619, n14620, n14621, n14622, n14623, n14624, n14625,
         n14626, n14627, n14628, n14629, n14630, n14631, n14632, n14633,
         n14634, n14635, n14636, n14637, n14638, n14639, n14640, n14641,
         n14642, n14643, n14644, n14645, n14646, n14647, n14648, n14649,
         n14650, n14651, n14652, n14653, n14654, n14655, n14656, n14657,
         n14658, n14659, n14660, n14661, n14662, n14663, n14664, n14665,
         n14666, n14667, n14668, n14669, n14670, n14671, n14672, n14673,
         n14674, n14675, n14676, n14677, n14678, n14679, n14680, n14681,
         n14682, n14683, n14684, n14685, n14686, n14687, n14688, n14689,
         n14690, n14691, n14692, n14693, n14694, n14695, n14696, n14697,
         n14698, n14699, n14700, n14701, n14702, n14703, n14704, n14705,
         n14706, n14707, n14708, n14709, n14710, n14711, n14712, n14713,
         n14714, n14715, n14716, n14717, n14718, n14719, n14720, n14721,
         n14722, n14723, n14724, n14725, n14726, n14727, n14728, n14729,
         n14730, n14731, n14732, n14733, n14734, n14735, n14736, n14737,
         n14738, n14739, n14740, n14741, n14742, n14743, n14744, n14745,
         n14746, n14747, n14748, n14749, n14750, n14751, n14752, n14753,
         n14754, n14755, n14756, n14757, n14758, n14759, n14760, n14761,
         n14762, n14763, n14764, n14765, n14766, n14767, n14768, n14769,
         n14770, n14771, n14772, n14773, n14774, n14775, n14776, n14777,
         n14778, n14779, n14780, n14781, n14782, n14783, n14784, n14785,
         n14786, n14787, n14788, n14789, n14790, n14791, n14792, n14793,
         n14794, n14795, n14796, n14797, n14798, n14799, n14800, n14801,
         n14802, n14803, n14804, n14805, n14806, n14807, n14808, n14809,
         n14810, n14811, n14812, n14813, n14814, n14815, n14816, n14817,
         n14818, n14819, n14820, n14821, n14822, n14823, n14824, n14825,
         n14826, n14827, n14828, n14829, n14830, n14831, n14832, n14833,
         n14834, n14835, n14836, n14837, n14838, n14839, n14840, n14841,
         n14842, n14843, n14844, n14845, n14846, n14847, n14848, n14849,
         n14850, n14851, n14852, n14853, n14854, n14855, n14856, n14857,
         n14858, n14859, n14860, n14861, n14862, n14863, n14864, n14865,
         n14866, n14867, n14868, n14869, n14870, n14871, n14872, n14873,
         n14874, n14875, n14876, n14877, n14878, n14879, n14880, n14881,
         n14882, n14883, n14884, n14885, n14886, n14887, n14888, n14889,
         n14890, n14891, n14892, n14893, n14894, n14895, n14896, n14897,
         n14898, n14899, n14900, n14901, n14902, n14903, n14904, n14905,
         n14906, n14907, n14908, n14909, n14910, n14911, n14912, n14913,
         n14914, n14915, n14916, n14917, n14918, n14919, n14920, n14921,
         n14922, n14923, n14924, n14925, n14926, n14927, n14928, n14929,
         n14930, n14931, n14932, n14933, n14934, n14935, n14936, n14937,
         n14938, n14939, n14940, n14941, n14942, n14943, n14944, n14945,
         n14946, n14947, n14948, n14949, n14950, n14951, n14952, n14953,
         n14954, n14955, n14956, n14957, n14958, n14959, n14960, n14961,
         n14962, n14963, n14964, n14965, n14966, n14967, n14968, n14969,
         n14970, n14971, n14972, n14973, n14974, n14975, n14976, n14977,
         n14978, n14979, n14980, n14981, n14982, n14983, n14984, n14985,
         n14986, n14987, n14988, n14989, n14990, n14991, n14992, n14993,
         n14994, n14995, n14996, n14997, n14998, n14999, n15000, n15001,
         n15002, n15003, n15004, n15005, n15006, n15007, n15008, n15009,
         n15010, n15011, n15012, n15013, n15014, n15015, n15016, n15017,
         n15018, n15019, n15020, n15021, n15022, n15023, n15024, n15025,
         n15026, n15027, n15028, n15029, n15030, n15031, n15032, n15033,
         n15034, n15035, n15036, n15037, n15038, n15039, n15040, n15041,
         n15042, n15043, n15044, n15045, n15046, n15047, n15048, n15049,
         n15050, n15051, n15052, n15053, n15054, n15055, n15056, n15057,
         n15058, n15059, n15060, n15061, n15062, n15063, n15064, n15065,
         n15066, n15067, n15068, n15069, n15070, n15071, n15072, n15073,
         n15074, n15075, n15076, n15077, n15078, n15079, n15080, n15081,
         n15082, n15083, n15084, n15085, n15086, n15087, n15088, n15089,
         n15090, n15091, n15092, n15093, n15094, n15095, n15096, n15097,
         n15098, n15099, n15100, n15101, n15102, n15103, n15104, n15105,
         n15106, n15107, n15108, n15109, n15110, n15111, n15112, n15113,
         n15114, n15115, n15116, n15117, n15118, n15119, n15120, n15121,
         n15122, n15123, n15124, n15125, n15126, n15127, n15128, n15129,
         n15130, n15131, n15132, n15133, n15134, n15135, n15136, n15137,
         n15138, n15139, n15140, n15141, n15142, n15143, n15144, n15145,
         n15146, n15147, n15148, n15149, n15150, n15151, n15152, n15153,
         n15154, n15155, n15156, n15157, n15158, n15159, n15160, n15161,
         n15162, n15163, n15164, n15165, n15166, n15167, n15168, n15169,
         n15170, n15171, n15172, n15173, n15174, n15175, n15176, n15177,
         n15178, n15179, n15180, n15181, n15182, n15183, n15184, n15185,
         n15186, n15187, n15188, n15189, n15190, n15191, n15192, n15193,
         n15194, n15195, n15196, n15197, n15198, n15199, n15200, n15201,
         n15202, n15203, n15204, n15205, n15206, n15207, n15208, n15209,
         n15210, n15211, n15212, n15213, n15214, n15215, n15216, n15217,
         n15218, n15219, n15220, n15221, n15222, n15223, n15224, n15225,
         n15226, n15227, n15228, n15229, n15230, n15231, n15232, n15233,
         n15234, n15235, n15236, n15237, n15238, n15239, n15240, n15241,
         n15242, n15243, n15244, n15245, n15246, n15247, n15248, n15249,
         n15250, n15251, n15252, n15253, n15254, n15255, n15256, n15257,
         n15258, n15259, n15260, n15261, n15262, n15263, n15264, n15265,
         n15266, n15267, n15268, n15269, n15270, n15271, n15272, n15273,
         n15274, n15275, n15276, n15277, n15278, n15279, n15280, n15281,
         n15282, n15283, n15284, n15285, n15286, n15287, n15288, n15289,
         n15290, n15291, n15292, n15293, n15294, n15295, n15296, n15297,
         n15298, n15299, n15300, n15301, n15302, n15303, n15304, n15305,
         n15306, n15307, n15308, n15309, n15310, n15311, n15312, n15313,
         n15314, n15315, n15316, n15317, n15318, n15319, n15320, n15321,
         n15322, n15323, n15324, n15325, n15326, n15327, n15328, n15329,
         n15330, n15331, n15332, n15333, n15334, n15335, n15336, n15337,
         n15338, n15339, n15340, n15341, n15342, n15343, n15344, n15345,
         n15346, n15347, n15348, n15349, n15350, n15351, n15352, n15353,
         n15354, n15355, n15356, n15357, n15358, n15359, n15360, n15361,
         n15362, n15363, n15364, n15365, n15366, n15367, n15368, n15369,
         n15370, n15371, n15372, n15373, n15374, n15375, n15376, n15377,
         n15378, n15379, n15380, n15381, n15382, n15383, n15384, n15385,
         n15386, n15387, n15388, n15389, n15390, n15391, n15392, n15393,
         n15394, n15395, n15396, n15397, n15398, n15399, n15400, n15401,
         n15402, n15403, n15404, n15405, n15406, n15407, n15408, n15409,
         n15410, n15411, n15412, n15413, n15414, n15415, n15416, n15417,
         n15418, n15419, n15420, n15421, n15422, n15423, n15424, n15425,
         n15426, n15427, n15428, n15429, n15430, n15431, n15432, n15433,
         n15434, n15435, n15436, n15437, n15438, n15439, n15440, n15441,
         n15442, n15443, n15444, n15445, n15446, n15447, n15448, n15449,
         n15450, n15451, n15452, n15453, n15454, n15455, n15456, n15457,
         n15458, n15459, n15460, n15461, n15462, n15463, n15464, n15465,
         n15466, n15467, n15468, n15469, n15470, n15471, n15472, n15473,
         n15474, n15475, n15476, n15477, n15478, n15479, n15480, n15481,
         n15482, n15483, n15484, n15485, n15486, n15487, n15488, n15489,
         n15490, n15491, n15492, n15493, n15494, n15495, n15496, n15497,
         n15498, n15499, n15500, n15501, n15502, n15503, n15504, n15505,
         n15506, n15507, n15508, n15509, n15510, n15511, n15512, n15513,
         n15514, n15515, n15516, n15517, n15518, n15519, n15520, n15521,
         n15522, n15523, n15524, n15525, n15526, n15527, n15528, n15529,
         n15530, n15531, n15532, n15533, n15534, n15535, n15536, n15537,
         n15538, n15539, n15540, n15541, n15542, n15543, n15544, n15545,
         n15546, n15547, n15548, n15549, n15550, n15551, n15552, n15553,
         n15554, n15555, n15556, n15557, n15558, n15559, n15560, n15561,
         n15562, n15563, n15564, n15565, n15566, n15567, n15568, n15569,
         n15570, n15571, n15572, n15573, n15574, n15575, n15576, n15577,
         n15578, n15579, n15580, n15581, n15582, n15583, n15584, n15585,
         n15586, n15587, n15588, n15589, n15590, n15591, n15592, n15593,
         n15594, n15595, n15596, n15597, n15598, n15599, n15600, n15601,
         n15602, n15603, n15604, n15605, n15606, n15607, n15608, n15609,
         n15610, n15611, n15612, n15613, n15614, n15615, n15616, n15617,
         n15618, n15619, n15620, n15621, n15622, n15623, n15624, n15625,
         n15626, n15627, n15628, n15629, n15630, n15631, n15632, n15633,
         n15634, n15635, n15636, n15637, n15638, n15639, n15640, n15641,
         n15642, n15643, n15644, n15645, n15646, n15647, n15648, n15649,
         n15650, n15651, n15652, n15653, n15654, n15655, n15656, n15657,
         n15658, n15659, n15660, n15661, n15662, n15663, n15664, n15665,
         n15666, n15667, n15668, n15669, n15670, n15671, n15672, n15673,
         n15674, n15675, n15676, n15677, n15678, n15679, n15680, n15681,
         n15682, n15683, n15684, n15685, n15686, n15687, n15688, n15689,
         n15690, n15691, n15692, n15693, n15694, n15695, n15696, n15697,
         n15698, n15699, n15700, n15701, n15702, n15703, n15704, n15705,
         n15706, n15707, n15708, n15709, n15710, n15711, n15712, n15713,
         n15714, n15715, n15716, n15717, n15718, n15719, n15720, n15721,
         n15722, n15723, n15724, n15725, n15726, n15727, n15728, n15729,
         n15730, n15731, n15732, n15733, n15734, n15735, n15736, n15737,
         n15738, n15739, n15740, n15741, n15742, n15743, n15744, n15745,
         n15746, n15747, n15748, n15749, n15750, n15751, n15752, n15753,
         n15754, n15755, n15756, n15757, n15758, n15759, n15760, n15761,
         n15762, n15763, n15764, n15765, n15766, n15767, n15768, n15769,
         n15770, n15771, n15772, n15773, n15774, n15775, n15776, n15777,
         n15778, n15779, n15780, n15781, n15782, n15783, n15784, n15785,
         n15786, n15787, n15788, n15789, n15790, n15791, n15792, n15793,
         n15794, n15795, n15796, n15797, n15798, n15799, n15800, n15801,
         n15802, n15803, n15804, n15805, n15806, n15807, n15808, n15809,
         n15810, n15811, n15812, n15813, n15814, n15815, n15816, n15817,
         n15818, n15819, n15820, n15821, n15822, n15823, n15824, n15825,
         n15826, n15827, n15828, n15829, n15830, n15831, n15832, n15833,
         n15834, n15835, n15836, n15837, n15838, n15839, n15840, n15841,
         n15842, n15843, n15844, n15845, n15846, n15847, n15848, n15849,
         n15850, n15851, n15852, n15853, n15854, n15855, n15856, n15857,
         n15858, n15859, n15860, n15861, n15862, n15863, n15864, n15865,
         n15866, n15867, n15868, n15869, n15870, n15871, n15872, n15873,
         n15874, n15875, n15876, n15877, n15878, n15879, n15880, n15881,
         n15882, n15883, n15884, n15885, n15886, n15887, n15888, n15889,
         n15890, n15891, n15892, n15893, n15894, n15895, n15896, n15897,
         n15898, n15899, n15900, n15901, n15902, n15903, n15904, n15905,
         n15906, n15907, n15908, n15909, n15910, n15911, n15912, n15913,
         n15914, n15915, n15916, n15917, n15918, n15919, n15920, n15921,
         n15922, n15923, n15924, n15925, n15926, n15927, n15928, n15929,
         n15930, n15931, n15932, n15933, n15934, n15935, n15936, n15937,
         n15938, n15939, n15940, n15941, n15942, n15943, n15944, n15945,
         n15946, n15947, n15948, n15949, n15950, n15951, n15952, n15953,
         n15954, n15955, n15956, n15957, n15958, n15959, n15960, n15961,
         n15962, n15963, n15964, n15965, n15966, n15967, n15968, n15969,
         n15970, n15971, n15972, n15973, n15974, n15975, n15976, n15977,
         n15978, n15979, n15980, n15981, n15982, n15983, n15984, n15985,
         n15986, n15987, n15988, n15989, n15990, n15991, n15992, n15993,
         n15994, n15995, n15996, n15997, n15998, n15999, n16000, n16001,
         n16002, n16003, n16004, n16005, n16006, n16007, n16008, n16009,
         n16010, n16011, n16012, n16013, n16014, n16015, n16016, n16017,
         n16018, n16019, n16020, n16021, n16022, n16023, n16024, n16025,
         n16026, n16027, n16028, n16029, n16030, n16031, n16032, n16033,
         n16034, n16035, n16036, n16037, n16038, n16039, n16040, n16041,
         n16042, n16043, n16044, n16045, n16046, n16047, n16048, n16049,
         n16050, n16051, n16052, n16053, n16054, n16055, n16056, n16057,
         n16058, n16059, n16060, n16061, n16062, n16063, n16064, n16065,
         n16066, n16067, n16068, n16069, n16070, n16071, n16072, n16073,
         n16074, n16075, n16076, n16077, n16078, n16079, n16080, n16081,
         n16082, n16083, n16084, n16085, n16086, n16087, n16088, n16089,
         n16090, n16091, n16092, n16093, n16094, n16095, n16096, n16097,
         n16098, n16099, n16100, n16101, n16102, n16103, n16104, n16105,
         n16106, n16107, n16108, n16109, n16110, n16111, n16112, n16113,
         n16114, n16115, n16116, n16117, n16118, n16119, n16120, n16121,
         n16122, n16123, n16124, n16125, n16126, n16127, n16128, n16129,
         n16130, n16131, n16132, n16133, n16134, n16135, n16136, n16137,
         n16138, n16139, n16140, n16141, n16142, n16143, n16144, n16145,
         n16146, n16147, n16148, n16149, n16150, n16151, n16152, n16153,
         n16154, n16155, n16156, n16157, n16158, n16159, n16160, n16161,
         n16162, n16163, n16164, n16165, n16166, n16167, n16168, n16169,
         n16170, n16171, n16172, n16173, n16174, n16175, n16176, n16177,
         n16178, n16179, n16180, n16181, n16182, n16183, n16184, n16185,
         n16186, n16187, n16188, n16189, n16190, n16191, n16192, n16193,
         n16194, n16195, n16196, n16197, n16198, n16199, n16200, n16201,
         n16202, n16203, n16204, n16205, n16206, n16207, n16208, n16209,
         n16210, n16211, n16212, n16213, n16214, n16215, n16216, n16217,
         n16218, n16219, n16220, n16221, n16222, n16223, n16224, n16225,
         n16226, n16227, n16228, n16229, n16230, n16231, n16232, n16233,
         n16234, n16235, n16236, n16237, n16238, n16239, n16240, n16241,
         n16242, n16243, n16244, n16245, n16246, n16247, n16248, n16249,
         n16250, n16251, n16252, n16253, n16254, n16255, n16256, n16257,
         n16258, n16259, n16260, n16261, n16262, n16263, n16264, n16265,
         n16266, n16267, n16268, n16269, n16270, n16271, n16272, n16273,
         n16274, n16275, n16276, n16277, n16278, n16279, n16280, n16281,
         n16282, n16283, n16284, n16285, n16286, n16287, n16288, n16289,
         n16290, n16291, n16292, n16293, n16294, n16295, n16296, n16297,
         n16298, n16299, n16300, n16301, n16302, n16303, n16304, n16305,
         n16306, n16307, n16308, n16309, n16310, n16311, n16312, n16313,
         n16314, n16315, n16316, n16317, n16318, n16319, n16320, n16321,
         n16322, n16323, n16324, n16325, n16326, n16327, n16328, n16329,
         n16330, n16331, n16332, n16333, n16334, n16335, n16336, n16337,
         n16338, n16339, n16340, n16341, n16342, n16343, n16344, n16345,
         n16346, n16347, n16348, n16349, n16350, n16351, n16352, n16353,
         n16354, n16355, n16356, n16357, n16358, n16359, n16360, n16361,
         n16362, n16363, n16364, n16365, n16366, n16367, n16368, n16369,
         n16370, n16371, n16372, n16373, n16374, n16375, n16376, n16377,
         n16378, n16379, n16380, n16381, n16382, n16383, n16384, n16385,
         n16386, n16387, n16388, n16389, n16390, n16391, n16392, n16393,
         n16394, n16395, n16396, n16397, n16398, n16399, n16400, n16401,
         n16402, n16403, n16404, n16405, n16406, n16407, n16408, n16409,
         n16410, n16411, n16412, n16413, n16414, n16415, n16416, n16417,
         n16418, n16419, n16420, n16421, n16422, n16423, n16424, n16425,
         n16426, n16427, n16428, n16429, n16430, n16431, n16432, n16433,
         n16434, n16435, n16436, n16437, n16438, n16439, n16440, n16441,
         n16442, n16443, n16444, n16445, n16446, n16447, n16448, n16449,
         n16450, n16451, n16452, n16453, n16454, n16455, n16456, n16457,
         n16458, n16459, n16460, n16461, n16462, n16463, n16464, n16465,
         n16466, n16467, n16468, n16469, n16470, n16471, n16472, n16473,
         n16474, n16475, n16476, n16477, n16478, n16479, n16480, n16481,
         n16482, n16483, n16484, n16485, n16486, n16487, n16488, n16489,
         n16490, n16491, n16492, n16493, n16494, n16495, n16496, n16497,
         n16498, n16499, n16500, n16501, n16502, n16503, n16504, n16505,
         n16506, n16507, n16508, n16509, n16510, n16511, n16512, n16513,
         n16514, n16515, n16516, n16517, n16518, n16519, n16520, n16521,
         n16522, n16523, n16524, n16525, n16526, n16527, n16528, n16529,
         n16530, n16531, n16532, n16533, n16534, n16535, n16536, n16537,
         n16538, n16539, n16540, n16541, n16542, n16543, n16544, n16545,
         n16546, n16547, n16548, n16549, n16550, n16551, n16552, n16553,
         n16554, n16555, n16556, n16557, n16558, n16559, n16560, n16561,
         n16562, n16563, n16564, n16565, n16566, n16567, n16568, n16569,
         n16570, n16571, n16572, n16573, n16574, n16575, n16576, n16577,
         n16578, n16579, n16580, n16581, n16582, n16583, n16584, n16585,
         n16586, n16587, n16588, n16589, n16590, n16591, n16592, n16593,
         n16594, n16595, n16596, n16597, n16598, n16599, n16600, n16601,
         n16602, n16603, n16604, n16605, n16606, n16607, n16608, n16609,
         n16610, n16611, n16612, n16613, n16614, n16615, n16616, n16617,
         n16618, n16619, n16620, n16621, n16622, n16623, n16624, n16625,
         n16626, n16627, n16628, n16629, n16630, n16631, n16632, n16633,
         n16634, n16635, n16636, n16637, n16638, n16639, n16640, n16641,
         n16642, n16643, n16644, n16645, n16646, n16647, n16648, n16649,
         n16650, n16651, n16652, n16653, n16654, n16655, n16656, n16657,
         n16658, n16659, n16660, n16661, n16662, n16663, n16664, n16665,
         n16666, n16667, n16668, n16669, n16670, n16671, n16672, n16673,
         n16674, n16675, n16676, n16677, n16678, n16679, n16680, n16681,
         n16682, n16683, n16684, n16685, n16686, n16687, n16688, n16689,
         n16690, n16691, n16692, n16693, n16694, n16695, n16696, n16697,
         n16698, n16699, n16700, n16701, n16702, n16703, n16704, n16705,
         n16706, n16707, n16708, n16709, n16710, n16711, n16712, n16713,
         n16714, n16715, n16716, n16717, n16718, n16719, n16720, n16721,
         n16722, n16723, n16724, n16725, n16726, n16727, n16728, n16729,
         n16730, n16731, n16732, n16733, n16734, n16735, n16736, n16737,
         n16738, n16739, n16740, n16741, n16742, n16743, n16744, n16745,
         n16746, n16747, n16748, n16749, n16750, n16751, n16752, n16753,
         n16754, n16755, n16756, n16757, n16758, n16759, n16760, n16761,
         n16762, n16763, n16764, n16765, n16766, n16767, n16768, n16769,
         n16770, n16771, n16772, n16773, n16774, n16775, n16776, n16777,
         n16778, n16779, n16780, n16781, n16782, n16783, n16784, n16785,
         n16786, n16787, n16788, n16789, n16790, n16791, n16792, n16793,
         n16794, n16795, n16796, n16797, n16798, n16799, n16800, n16801,
         n16802, n16803, n16804, n16805, n16806, n16807, n16808, n16809,
         n16810, n16811, n16812, n16813, n16814, n16815, n16816, n16817,
         n16818, n16819, n16820, n16821, n16822, n16823, n16824, n16825,
         n16826, n16827, n16828, n16829, n16830, n16831, n16832, n16833,
         n16834, n16835, n16836, n16837, n16838, n16839, n16840, n16841,
         n16842, n16843, n16844, n16845, n16846, n16847, n16848, n16849,
         n16850, n16851, n16852, n16853, n16854, n16855, n16856, n16857,
         n16858, n16859, n16860, n16861, n16862, n16863, n16864, n16865,
         n16866, n16867, n16868, n16869, n16870, n16871, n16872, n16873,
         n16874, n16875, n16876, n16877, n16878, n16879, n16880, n16881,
         n16882, n16883, n16884, n16885, n16886, n16887, n16888, n16889,
         n16890, n16891, n16892, n16893, n16894, n16895, n16896, n16897,
         n16898, n16899, n16900, n16901, n16902, n16903, n16904, n16905,
         n16906, n16907, n16908, n16909, n16910, n16911, n16912, n16913,
         n16914, n16915, n16916, n16917, n16918, n16919, n16920, n16921,
         n16922, n16923, n16924, n16925, n16926, n16927, n16928, n16929,
         n16930, n16931, n16932, n16933, n16934, n16935, n16936, n16937,
         n16938, n16939, n16940, n16941, n16942, n16943, n16944, n16945,
         n16946, n16947, n16948, n16949, n16950, n16951, n16952, n16953,
         n16954, n16955, n16956, n16957, n16958, n16959, n16960, n16961,
         n16962, n16963, n16964, n16965, n16966, n16967, n16968, n16969,
         n16970, n16971, n16972, n16973, n16974, n16975, n16976, n16977,
         n16978, n16979, n16980, n16981, n16982, n16983, n16984, n16985,
         n16986, n16987, n16988, n16989, n16990, n16991, n16992, n16993,
         n16994, n16995, n16996, n16997, n16998, n16999, n17000, n17001,
         n17002, n17003, n17004, n17005, n17006, n17007, n17008, n17009,
         n17010, n17011, n17012, n17013, n17014, n17015, n17016, n17017,
         n17018, n17019, n17020, n17021, n17022, n17023, n17024, n17025,
         n17026, n17027, n17028, n17029, n17030, n17031, n17032, n17033,
         n17034, n17035, n17036, n17037, n17038, n17039, n17040, n17041,
         n17042, n17043, n17044, n17045, n17046, n17047, n17048, n17049,
         n17050, n17051, n17052, n17053, n17054, n17055, n17056, n17057,
         n17058, n17059, n17060, n17061, n17062, n17063, n17064, n17065,
         n17066, n17067, n17068, n17069, n17070, n17071, n17072, n17073,
         n17074, n17075, n17076, n17077, n17078, n17079, n17080, n17081,
         n17082, n17083, n17084, n17085, n17086, n17087, n17088, n17089,
         n17090, n17091, n17092, n17093, n17094, n17095, n17096, n17097,
         n17098, n17099, n17100, n17101, n17102, n17103, n17104, n17105,
         n17106, n17107, n17108, n17109, n17110, n17111, n17112, n17113,
         n17114, n17115, n17116, n17117, n17118, n17119, n17120, n17121,
         n17122, n17123, n17124, n17125, n17126, n17127, n17128, n17129,
         n17130, n17131, n17132, n17133, n17134, n17135, n17136, n17137,
         n17138, n17139, n17140, n17141, n17142, n17143, n17144, n17145,
         n17146, n17147, n17148, n17149, n17150, n17151, n17152, n17153,
         n17154, n17155, n17156, n17157, n17158, n17159, n17160, n17161,
         n17162, n17163, n17164, n17165, n17166, n17167, n17168, n17169,
         n17170, n17171, n17172, n17173, n17174, n17175, n17176, n17177,
         n17178, n17179, n17180, n17181, n17182, n17183, n17184, n17185,
         n17186, n17187, n17188, n17189, n17190, n17191, n17192, n17193,
         n17194, n17195, n17196, n17197, n17198, n17199, n17200, n17201,
         n17202, n17203, n17204, n17205, n17206, n17207, n17208, n17209,
         n17210, n17211, n17212, n17213, n17214, n17215, n17216, n17217,
         n17218, n17219, n17220, n17221, n17222, n17223, n17224, n17225,
         n17226, n17227, n17228, n17229, n17230, n17231, n17232, n17233,
         n17234, n17235, n17236, n17237, n17238, n17239, n17240, n17241,
         n17242, n17243, n17244, n17245, n17246, n17247, n17248, n17249,
         n17250, n17251, n17252, n17253, n17254, n17255, n17256, n17257,
         n17258, n17259, n17260, n17261, n17262, n17263, n17264, n17265,
         n17266, n17267, n17268, n17269, n17270, n17271, n17272, n17273,
         n17274, n17275, n17276, n17277, n17278, n17279, n17280, n17281,
         n17282, n17283, n17284, n17285, n17286, n17287, n17288, n17289,
         n17290, n17291, n17292, n17293, n17294, n17295, n17296, n17297,
         n17298, n17299, n17300, n17301, n17302, n17303, n17304, n17305,
         n17306, n17307, n17308, n17309, n17310, n17311, n17312, n17313,
         n17314, n17315, n17316, n17317, n17318, n17319, n17320, n17321,
         n17322, n17323, n17324, n17325, n17326, n17327, n17328, n17329,
         n17330, n17331, n17332, n17333, n17334, n17335, n17336, n17337,
         n17338, n17339, n17340, n17341, n17342, n17343, n17344, n17345,
         n17346, n17347, n17348, n17349, n17350, n17351, n17352, n17353,
         n17354, n17355, n17356, n17357, n17358, n17359, n17360, n17361,
         n17362, n17363, n17364, n17365, n17366, n17367, n17368, n17369,
         n17370, n17371, n17372, n17373, n17374, n17375, n17376, n17377,
         n17378, n17379, n17380, n17381, n17382, n17383, n17384, n17385,
         n17386, n17387, n17388, n17389, n17390, n17391, n17392, n17393,
         n17394, n17395, n17396, n17397, n17398, n17399, n17400, n17401,
         n17402, n17403, n17404, n17405, n17406, n17407, n17408, n17409,
         n17410, n17411, n17412, n17413, n17414, n17415, n17416, n17417,
         n17418, n17419, n17420, n17421, n17422, n17423, n17424, n17425,
         n17426, n17427, n17428, n17429, n17430, n17431, n17432, n17433,
         n17434, n17435, n17436, n17437, n17438, n17439, n17440, n17441,
         n17442, n17443, n17444, n17445, n17446, n17447, n17448, n17449,
         n17450, n17451, n17452, n17453, n17454, n17455, n17456, n17457,
         n17458, n17459, n17460, n17461, n17462, n17463, n17464, n17465,
         n17466, n17467, n17468, n17469, n17470, n17471, n17472, n17473,
         n17474, n17475, n17476, n17477, n17478, n17479, n17480, n17481,
         n17482, n17483, n17484, n17485, n17486, n17487, n17488, n17489,
         n17490, n17491, n17492, n17493, n17494, n17495, n17496, n17497,
         n17498, n17499, n17500, n17501, n17502, n17503, n17504, n17505,
         n17506, n17507, n17508, n17509, n17510, n17511, n17512, n17513,
         n17514, n17515, n17516, n17517, n17518, n17519, n17520, n17521,
         n17522, n17523, n17524, n17525, n17526, n17527, n17528, n17529,
         n17530, n17531, n17532, n17533, n17534, n17535, n17536, n17537,
         n17538, n17539, n17540, n17541, n17542, n17543, n17544, n17545,
         n17546, n17547, n17548, n17549, n17550, n17551, n17552, n17553,
         n17554, n17555, n17556, n17557, n17558, n17559, n17560, n17561,
         n17562, n17563, n17564, n17565, n17566, n17567, n17568, n17569,
         n17570, n17571, n17572, n17573, n17574, n17575, n17576, n17577,
         n17578, n17579, n17580, n17581, n17582, n17583, n17584, n17585,
         n17586, n17587, n17588, n17589, n17590, n17591, n17592, n17593,
         n17594, n17595, n17596, n17597, n17598, n17599, n17600, n17601,
         n17602, n17603, n17604, n17605, n17606, n17607, n17608, n17609,
         n17610, n17611, n17612, n17613, n17614, n17615, n17616, n17617,
         n17618, n17619, n17620, n17621, n17622, n17623, n17624, n17625,
         n17626, n17627, n17628, n17629, n17630, n17631, n17632, n17633,
         n17634, n17635, n17636, n17637, n17638, n17639, n17640, n17641,
         n17642, n17643, n17644, n17645, n17646, n17647, n17648, n17649,
         n17650, n17651, n17652, n17653, n17654, n17655, n17656, n17657,
         n17658, n17659, n17660, n17661, n17662, n17663, n17664, n17665,
         n17666, n17667, n17668, n17669, n17670, n17671, n17672, n17673,
         n17674, n17675, n17676, n17677, n17678, n17679, n17680, n17681,
         n17682, n17683, n17684, n17685, n17686, n17687, n17688, n17689,
         n17690, n17691, n17692, n17693, n17694, n17695, n17696, n17697,
         n17698, n17699, n17700, n17701, n17702, n17703, n17704, n17705,
         n17706, n17707, n17708, n17709, n17710, n17711, n17712, n17713,
         n17714, n17715, n17716, n17717, n17718, n17719, n17720, n17721,
         n17722, n17723, n17724, n17725, n17726, n17727, n17728, n17729,
         n17730, n17731, n17732, n17733, n17734, n17735, n17736, n17737,
         n17738, n17739, n17740, n17741, n17742, n17743, n17744, n17745,
         n17746, n17747, n17748, n17749, n17750, n17751, n17752, n17753,
         n17754, n17755, n17756, n17757, n17758, n17759, n17760, n17761,
         n17762, n17763, n17764, n17765, n17766, n17767, n17768, n17769,
         n17770, n17771, n17772, n17773, n17774, n17775, n17776, n17777,
         n17778, n17779, n17780, n17781, n17782, n17783, n17784, n17785,
         n17786, n17787, n17788, n17789, n17790, n17791, n17792, n17793,
         n17794, n17795, n17796, n17797, n17798, n17799, n17800, n17801,
         n17802, n17803, n17804, n17805, n17806, n17807, n17808, n17809,
         n17810, n17811, n17812, n17813, n17814, n17815, n17816, n17817,
         n17818, n17819, n17820, n17821, n17822, n17823, n17824, n17825,
         n17826, n17827, n17828, n17829, n17830, n17831, n17832, n17833,
         n17834, n17835, n17836, n17837, n17838, n17839, n17840, n17841,
         n17842, n17843, n17844, n17845, n17846, n17847, n17848, n17849,
         n17850, n17851, n17852, n17853, n17854, n17855, n17856, n17857,
         n17858, n17859, n17860, n17861, n17862, n17863, n17864, n17865,
         n17866, n17867, n17868, n17869, n17870, n17871, n17872, n17873,
         n17874, n17875, n17876, n17877, n17878, n17879, n17880, n17881,
         n17882, n17883, n17884, n17885, n17886, n17887, n17888, n17889,
         n17890, n17891, n17892, n17893, n17894, n17895, n17896, n17897,
         n17898, n17899, n17900, n17901, n17902, n17903, n17904, n17905,
         n17906, n17907, n17908, n17909, n17910, n17911, n17912, n17913,
         n17914, n17915, n17916, n17917, n17918, n17919, n17920, n17921,
         n17922, n17923, n17924, n17925, n17926, n17927, n17928, n17929,
         n17930, n17931, n17932, n17933, n17934, n17935, n17936, n17937,
         n17938, n17939, n17940, n17941, n17942, n17943, n17944, n17945,
         n17946, n17947, n17948, n17949, n17950, n17951, n17952, n17953,
         n17954, n17955, n17956, n17957, n17958, n17959, n17960, n17961,
         n17962, n17963, n17964, n17965, n17966, n17967, n17968, n17969,
         n17970, n17971, n17972, n17973, n17974, n17975, n17976, n17977,
         n17978, n17979, n17980, n17981, n17982, n17983, n17984, n17985,
         n17986, n17987, n17988, n17989, n17990, n17991, n17992, n17993,
         n17994, n17995, n17996, n17997, n17998, n17999, n18000, n18001,
         n18002, n18003, n18004, n18005, n18006, n18007, n18008, n18009,
         n18010, n18011, n18012, n18013, n18014, n18015, n18016, n18017,
         n18018, n18019, n18020, n18021, n18022, n18023, n18024, n18025,
         n18026, n18027, n18028, n18029, n18030, n18031, n18032, n18033,
         n18034, n18035, n18036, n18037, n18038, n18039, n18040, n18041,
         n18042, n18043, n18044, n18045, n18046, n18047, n18048, n18049,
         n18050, n18051, n18052, n18053, n18054, n18055, n18056, n18057,
         n18058, n18059, n18060, n18061, n18062, n18063, n18064, n18065,
         n18066, n18067, n18068, n18069, n18070, n18071, n18072, n18073,
         n18074, n18075, n18076, n18077, n18078, n18079, n18080, n18081,
         n18082, n18083, n18084, n18085, n18086, n18087, n18088, n18089,
         n18090, n18091, n18092, n18093, n18094, n18095, n18096, n18097,
         n18098, n18099, n18100, n18101, n18102, n18103, n18104, n18105,
         n18106, n18107, n18108, n18109, n18110, n18111, n18112, n18113,
         n18114, n18115, n18116, n18117, n18118, n18119, n18120, n18121,
         n18122, n18123, n18124, n18125, n18126, n18127, n18128, n18129,
         n18130, n18131, n18132, n18133, n18134, n18135, n18136, n18137,
         n18138, n18139, n18140, n18141, n18142, n18143, n18144, n18145,
         n18146, n18147, n18148, n18149, n18150, n18151, n18152, n18153,
         n18154, n18155, n18156, n18157, n18158, n18159, n18160, n18161,
         n18162, n18163, n18164, n18165, n18166, n18167, n18168, n18169,
         n18170, n18171, n18172, n18173, n18174, n18175, n18176, n18177,
         n18178, n18179, n18180, n18181, n18182, n18183, n18184, n18185,
         n18186, n18187, n18188, n18189, n18190, n18191, n18192, n18193,
         n18194, n18195, n18196, n18197, n18198, n18199, n18200, n18201,
         n18202, n18203, n18204, n18205, n18206, n18207, n18208, n18209,
         n18210, n18211, n18212, n18213, n18214, n18215, n18216, n18217,
         n18218, n18219, n18220, n18221, n18222, n18223, n18224, n18225,
         n18226, n18227, n18228, n18229, n18230, n18231, n18232, n18233,
         n18234, n18235, n18236, n18237, n18238, n18239, n18240, n18241,
         n18242, n18243, n18244, n18245, n18246, n18247, n18248, n18249,
         n18250, n18251, n18252, n18253, n18254, n18255, n18256, n18257,
         n18258, n18259, n18260, n18261, n18262, n18263, n18264, n18265,
         n18266, n18267, n18268, n18269, n18270, n18271, n18272, n18273,
         n18274, n18275, n18276, n18277, n18278, n18279, n18280, n18281,
         n18282, n18283, n18284, n18285, n18286, n18287, n18288, n18289,
         n18290, n18291, n18292, n18293, n18294, n18295, n18296, n18297,
         n18298, n18299, n18300, n18301, n18302, n18303, n18304, n18305,
         n18306, n18307, n18308, n18309, n18310, n18311, n18312, n18313,
         n18314, n18315, n18316, n18317, n18318, n18319, n18320, n18321,
         n18322, n18323, n18324, n18325, n18326, n18327, n18328, n18329,
         n18330, n18331, n18332, n18333, n18334, n18335, n18336, n18337,
         n18338, n18339, n18340, n18341, n18342, n18343, n18344, n18345,
         n18346, n18347, n18348, n18349, n18350, n18351, n18352, n18353,
         n18354, n18355, n18356, n18357, n18358, n18359, n18360, n18361,
         n18362, n18363, n18364, n18365, n18366, n18367, n18368, n18369,
         n18370, n18371, n18372, n18373, n18374, n18375, n18376, n18377,
         n18378, n18379, n18380, n18381, n18382, n18383, n18384, n18385,
         n18386, n18387, n18388, n18389, n18390, n18391, n18392, n18393,
         n18394, n18395, n18396, n18397, n18398, n18399, n18400, n18401,
         n18402, n18403, n18404, n18405, n18406, n18407, n18408, n18409,
         n18410, n18411, n18412, n18413, n18414, n18415, n18416, n18417,
         n18418, n18419, n18420, n18421, n18422, n18423, n18424, n18425,
         n18426, n18427, n18428, n18429, n18430, n18431, n18432, n18433,
         n18434, n18435, n18436, n18437, n18438, n18439, n18440, n18441,
         n18442, n18443, n18444, n18445, n18446, n18447, n18448, n18449,
         n18450, n18451, n18452, n18453, n18454, n18455, n18456, n18457,
         n18458, n18459, n18460, n18461, n18462, n18463, n18464, n18465,
         n18466, n18467, n18468, n18469, n18470, n18471, n18472, n18473,
         n18474, n18475, n18476, n18477, n18478, n18479, n18480, n18481,
         n18482, n18483, n18484, n18485, n18486, n18487, n18488, n18489,
         n18490, n18491, n18492, n18493, n18494, n18495, n18496, n18497,
         n18498, n18499, n18500, n18501, n18502, n18503, n18504, n18505,
         n18506, n18507, n18508, n18509, n18510, n18511, n18512, n18513,
         n18514, n18515, n18516, n18517, n18518, n18519, n18520, n18521,
         n18522, n18523, n18524, n18525, n18526, n18527, n18528, n18529,
         n18530, n18531, n18532, n18533, n18534, n18535, n18536, n18537,
         n18538, n18539, n18540, n18541, n18542, n18543, n18544, n18545,
         n18546, n18547, n18548, n18549, n18550, n18551, n18552, n18553,
         n18554, n18555, n18556, n18557, n18558, n18559, n18560, n18561,
         n18562, n18563, n18564, n18565, n18566, n18567, n18568, n18569,
         n18570, n18571, n18572, n18573, n18574, n18575, n18576, n18577,
         n18578, n18579, n18580, n18581, n18582, n18583, n18584, n18585,
         n18586, n18587, n18588, n18589, n18590, n18591, n18592, n18593,
         n18594, n18595, n18596, n18597, n18598, n18599, n18600, n18601,
         n18602, n18603, n18604, n18605, n18606, n18607, n18608, n18609,
         n18610, n18611, n18612, n18613, n18614, n18615, n18616, n18617,
         n18618, n18619, n18620, n18621, n18622, n18623, n18624, n18625,
         n18626, n18627, n18628, n18629, n18630, n18631, n18632, n18633,
         n18634, n18635, n18636, n18637, n18638, n18639, n18640, n18641,
         n18642, n18643, n18644, n18645, n18646, n18647, n18648, n18649,
         n18650, n18651, n18652, n18653, n18654, n18655, n18656, n18657,
         n18658, n18659, n18660, n18661, n18662, n18663, n18664, n18665,
         n18666, n18667, n18668, n18669, n18670, n18671, n18672, n18673,
         n18674, n18675, n18676, n18677, n18678, n18679, n18680, n18681,
         n18682, n18683, n18684, n18685, n18686, n18687, n18688, n18689,
         n18690, n18691, n18692, n18693, n18694, n18695, n18696, n18697,
         n18698, n18699, n18700, n18701, n18702, n18703, n18704, n18705,
         n18706, n18707, n18708, n18709, n18710, n18711, n18712, n18713,
         n18714, n18715, n18716, n18717, n18718, n18719, n18720, n18721,
         n18722, n18723, n18724, n18725, n18726, n18727, n18728, n18729,
         n18730, n18731, n18732, n18733, n18734, n18735, n18736, n18737,
         n18738, n18739, n18740, n18741, n18742, n18743, n18744, n18745,
         n18746, n18747, n18748, n18749, n18750, n18751, n18752, n18753,
         n18754, n18755, n18756, n18757, n18758, n18759, n18760, n18761,
         n18762, n18763, n18764, n18765, n18766, n18767, n18768, n18769,
         n18770, n18771, n18772, n18773, n18774, n18775, n18776, n18777,
         n18778, n18779, n18780, n18781, n18782, n18783, n18784, n18785,
         n18786, n18787, n18788, n18789, n18790, n18791, n18792, n18793,
         n18794, n18795, n18796, n18797, n18798, n18799, n18800, n18801,
         n18802, n18803, n18804, n18805, n18806, n18807, n18808, n18809,
         n18810, n18811, n18812, n18813, n18814, n18815, n18816, n18817,
         n18818, n18819, n18820, n18821, n18822, n18823, n18824, n18825,
         n18826, n18827, n18828, n18829, n18830, n18831, n18832, n18833,
         n18834, n18835, n18836, n18837, n18838, n18839, n18840, n18841,
         n18842, n18843, n18844, n18845, n18846, n18847, n18848, n18849,
         n18850, n18851, n18852, n18853, n18854, n18855, n18856, n18857,
         n18858, n18859, n18860, n18861, n18862, n18863, n18864, n18865,
         n18866, n18867, n18868, n18869, n18870, n18871, n18872, n18873,
         n18874, n18875, n18876, n18877, n18878, n18879, n18880, n18881,
         n18882, n18883, n18884, n18885, n18886, n18887, n18888, n18889,
         n18890, n18891, n18892, n18893, n18894, n18895, n18896, n18897,
         n18898, n18899, n18900, n18901, n18902, n18903, n18904, n18905,
         n18906, n18907, n18908, n18909, n18910, n18911, n18912, n18913,
         n18914, n18915, n18916, n18917, n18918, n18919, n18920, n18921,
         n18922, n18923, n18924, n18925, n18926, n18927, n18928, n18929,
         n18930, n18931, n18932, n18933, n18934, n18935, n18936, n18937,
         n18938, n18939, n18940, n18941, n18942, n18943, n18944, n18945,
         n18946, n18947, n18948, n18949, n18950, n18951, n18952, n18953,
         n18954, n18955, n18956, n18957, n18958, n18959, n18960, n18961,
         n18962, n18963, n18964, n18965, n18966, n18967, n18968, n18969,
         n18970, n18971, n18972, n18973, n18974, n18975, n18976, n18977,
         n18978, n18979, n18980, n18981, n18982, n18983, n18984, n18985,
         n18986, n18987, n18988, n18989, n18990, n18991, n18992, n18993,
         n18994, n18995, n18996, n18997, n18998, n18999, n19000, n19001,
         n19002, n19003, n19004, n19005, n19006, n19007, n19008, n19009,
         n19010, n19011, n19012, n19013, n19014, n19015, n19016, n19017,
         n19018, n19019, n19020, n19021, n19022, n19023, n19024, n19025,
         n19026, n19027, n19028, n19029, n19030, n19031, n19032, n19033,
         n19034, n19035, n19036, n19037, n19038, n19039, n19040, n19041,
         n19042, n19043, n19044, n19045, n19046, n19047, n19048, n19049,
         n19050, n19051, n19052, n19053, n19054, n19055, n19056, n19057,
         n19058, n19059, n19060, n19061, n19062, n19063, n19064, n19065,
         n19066, n19067, n19068, n19069, n19070, n19071, n19072, n19073,
         n19074, n19075, n19076, n19077, n19078, n19079, n19080, n19081,
         n19082, n19083, n19084, n19085, n19086, n19087, n19088, n19089,
         n19090, n19091, n19092, n19093, n19094, n19095, n19096, n19097,
         n19098, n19099, n19100, n19101, n19102, n19103, n19104, n19105,
         n19106, n19107, n19108, n19109, n19110, n19111, n19112, n19113,
         n19114, n19115, n19116, n19117, n19118, n19119, n19120, n19121,
         n19122, n19123, n19124, n19125, n19126, n19127, n19128, n19129,
         n19130, n19131, n19132, n19133, n19134, n19135, n19136, n19137,
         n19138, n19139, n19140, n19141, n19142, n19143, n19144, n19145,
         n19146, n19147, n19148, n19149, n19150, n19151, n19152, n19153,
         n19154, n19155, n19156, n19157, n19158, n19159, n19160, n19161,
         n19162, n19163, n19164, n19165, n19166, n19167, n19168, n19169,
         n19170, n19171, n19172, n19173, n19174, n19175, n19176, n19177,
         n19178, n19179, n19180, n19181, n19182, n19183, n19184, n19185,
         n19186, n19187, n19188, n19189, n19190, n19191, n19192, n19193,
         n19194, n19195, n19196, n19197, n19198, n19199, n19200, n19201,
         n19202, n19203, n19204, n19205, n19206, n19207, n19208, n19209,
         n19210, n19211, n19212, n19213, n19214, n19215, n19216, n19217,
         n19218, n19219, n19220, n19221, n19222, n19223, n19224, n19225,
         n19226, n19227, n19228, n19229, n19230, n19231, n19232, n19233,
         n19234, n19235, n19236, n19237, n19238, n19239, n19240, n19241,
         n19242, n19243, n19244, n19245, n19246, n19247, n19248, n19249,
         n19250, n19251, n19252, n19253, n19254, n19255, n19256, n19257,
         n19258, n19259, n19260, n19261, n19262, n19263, n19264, n19265,
         n19266, n19267, n19268, n19269, n19270, n19271, n19272, n19273,
         n19274, n19275, n19276, n19277, n19278, n19279, n19280, n19281,
         n19282, n19283, n19284, n19285, n19286, n19287, n19288, n19289,
         n19290, n19291, n19292, n19293, n19294, n19295, n19296, n19297,
         n19298, n19299, n19300, n19301, n19302, n19303, n19304, n19305,
         n19306, n19307, n19308, n19309, n19310, n19311, n19312, n19313,
         n19314, n19315, n19316, n19317, n19318, n19319, n19320, n19321,
         n19322, n19323, n19324, n19325, n19326, n19327, n19328, n19329,
         n19330, n19331, n19332, n19333, n19334, n19335, n19336, n19337,
         n19338, n19339, n19340, n19341, n19342, n19343, n19344, n19345,
         n19346, n19347, n19348, n19349, n19350, n19351, n19352, n19353,
         n19354, n19355, n19356, n19357, n19358, n19359, n19360, n19361,
         n19362, n19363, n19364, n19365, n19366, n19367, n19368, n19369,
         n19370, n19371, n19372, n19373, n19374, n19375, n19376, n19377,
         n19378, n19379, n19380, n19381, n19382, n19383, n19384, n19385,
         n19386, n19387, n19388, n19389, n19390, n19391, n19392, n19393,
         n19394, n19395, n19396, n19397, n19398, n19399, n19400, n19401,
         n19402, n19403, n19404, n19405, n19406, n19407, n19408, n19409,
         n19410, n19411, n19412, n19413, n19414, n19415, n19416, n19417,
         n19418, n19419, n19420, n19421, n19422, n19423, n19424, n19425,
         n19426, n19427, n19428, n19429, n19430, n19431, n19432, n19433,
         n19434, n19435, n19436, n19437, n19438, n19439, n19440, n19441,
         n19442, n19443, n19444, n19445, n19446, n19447, n19448, n19449,
         n19450, n19451, n19452, n19453, n19454, n19455, n19456, n19457,
         n19458, n19459, n19460, n19461, n19462, n19463, n19464, n19465,
         n19466, n19467, n19468, n19469, n19470, n19471, n19472, n19473,
         n19474, n19475, n19476, n19477, n19478, n19479, n19480, n19481,
         n19482, n19483, n19484, n19485, n19486, n19487, n19488, n19489,
         n19490, n19491, n19492, n19493, n19494, n19495, n19496, n19497,
         n19498, n19499, n19500, n19501, n19502, n19503, n19504, n19505,
         n19506, n19507, n19508, n19509, n19510, n19511, n19512, n19513,
         n19514, n19515, n19516, n19517, n19518, n19519, n19520, n19521,
         n19522, n19523, n19524, n19525, n19526, n19527, n19528, n19529,
         n19530, n19531, n19532, n19533, n19534, n19535, n19536, n19537,
         n19538, n19539, n19540, n19541, n19542, n19543, n19544, n19545,
         n19546, n19547, n19548, n19549, n19550, n19551, n19552, n19553,
         n19554, n19555, n19556, n19557, n19558, n19559, n19560, n19561,
         n19562, n19563, n19564, n19565, n19566, n19567, n19568, n19569,
         n19570, n19571, n19572, n19573, n19574, n19575, n19576, n19577,
         n19578, n19579, n19580, n19581, n19582, n19583, n19584, n19585,
         n19586, n19587, n19588, n19589, n19590, n19591, n19592, n19593,
         n19594, n19595, n19596, n19597, n19598, n19599, n19600, n19601,
         n19602, n19603, n19604, n19605, n19606, n19607, n19608, n19609,
         n19610, n19611, n19612, n19613, n19614, n19615, n19616, n19617,
         n19618, n19619, n19620, n19621, n19622, n19623, n19624, n19625,
         n19626, n19627, n19628, n19629, n19630, n19631, n19632, n19633,
         n19634, n19635, n19636, n19637, n19638, n19639, n19640, n19641,
         n19642, n19643, n19644, n19645, n19646, n19647, n19648, n19649,
         n19650, n19651, n19652, n19653, n19654, n19655, n19656, n19657,
         n19658, n19659, n19660, n19661, n19662, n19663, n19664, n19665,
         n19666, n19667, n19668, n19669, n19670, n19671, n19672, n19673,
         n19674, n19675, n19676, n19677, n19678, n19679, n19680, n19681,
         n19682, n19683, n19684, n19685, n19686, n19687, n19688, n19689,
         n19690, n19691, n19692, n19693, n19694, n19695, n19696, n19697,
         n19698, n19699, n19700, n19701, n19702, n19703, n19704, n19705,
         n19706, n19707, n19708, n19709, n19710, n19711, n19712, n19713,
         n19714, n19715, n19716, n19717, n19718, n19719, n19720, n19721,
         n19722, n19723, n19724, n19725, n19726, n19727, n19728, n19729,
         n19730, n19731, n19732, n19733, n19734, n19735, n19736, n19737,
         n19738, n19739, n19740, n19741, n19742, n19743, n19744, n19745,
         n19746, n19747, n19748, n19749, n19750, n19751, n19752, n19753,
         n19754, n19755, n19756, n19757, n19758, n19759, n19760, n19761,
         n19762, n19763, n19764, n19765, n19766, n19767, n19768, n19769,
         n19770, n19771, n19772, n19773, n19774, n19775, n19776, n19777,
         n19778, n19779, n19780, n19781, n19782, n19783, n19784, n19785,
         n19786, n19787, n19788, n19789, n19790, n19791, n19792, n19793,
         n19794, n19795, n19796, n19797, n19798, n19799, n19800, n19801,
         n19802, n19803, n19804, n19805, n19806, n19807, n19808, n19809,
         n19810, n19811, n19812, n19813, n19814, n19815, n19816, n19817,
         n19818, n19819, n19820, n19821, n19822, n19823, n19824, n19825,
         n19826, n19827, n19828, n19829, n19830, n19831, n19832, n19833,
         n19834, n19835, n19836, n19837, n19838, n19839, n19840, n19841,
         n19842, n19843, n19844, n19845, n19846, n19847, n19848, n19849,
         n19850, n19851, n19852, n19853, n19854, n19855, n19856, n19857,
         n19858, n19859, n19860, n19861, n19862, n19863, n19864, n19865,
         n19866, n19867, n19868, n19869, n19870, n19871, n19872, n19873,
         n19874, n19875, n19876, n19877, n19878, n19879, n19880, n19881,
         n19882, n19883, n19884, n19885, n19886, n19887, n19888, n19889,
         n19890, n19891, n19892, n19893, n19894, n19895, n19896, n19897,
         n19898, n19899, n19900, n19901, n19902, n19903, n19904, n19905,
         n19906, n19907, n19908, n19909, n19910, n19911, n19912, n19913,
         n19914, n19915, n19916, n19917, n19918, n19919, n19920, n19921,
         n19922, n19923, n19924, n19925, n19926, n19927, n19928, n19929,
         n19930, n19931, n19932, n19933, n19934, n19935, n19936, n19937,
         n19938, n19939, n19940, n19941, n19942, n19943, n19944, n19945,
         n19946, n19947, n19948, n19949, n19950, n19951, n19952, n19953,
         n19954, n19955, n19956, n19957, n19958, n19959, n19960, n19961,
         n19962, n19963, n19964, n19965, n19966, n19967, n19968, n19969,
         n19970, n19971, n19972, n19973, n19974, n19975, n19976, n19977,
         n19978, n19979, n19980, n19981, n19982, n19983, n19984, n19985,
         n19986, n19987, n19988, n19989, n19990, n19991, n19992, n19993,
         n19994, n19995, n19996, n19997, n19998, n19999, n20000, n20001,
         n20002, n20003, n20004, n20005, n20006, n20007, n20008, n20009,
         n20010, n20011, n20012, n20013, n20014, n20015, n20016, n20017,
         n20018, n20019, n20020, n20021, n20022, n20023, n20024, n20025,
         n20026, n20027, n20028, n20029, n20030, n20031, n20032, n20033,
         n20034, n20035, n20036, n20037, n20038, n20039, n20040, n20041,
         n20042, n20043, n20044, n20045, n20046, n20047, n20048, n20049,
         n20050, n20051, n20052, n20053, n20054, n20055, n20056, n20057,
         n20058, n20059, n20060, n20061, n20062, n20063, n20064, n20065,
         n20066, n20067, n20068, n20069, n20070, n20071, n20072, n20073,
         n20074, n20075, n20076, n20077, n20078, n20079, n20080, n20081,
         n20082, n20083, n20084, n20085, n20086, n20087, n20088, n20089,
         n20090, n20091, n20092, n20093, n20094, n20095, n20096, n20097,
         n20098, n20099, n20100, n20101, n20102, n20103, n20104, n20105,
         n20106, n20107, n20108, n20109, n20110, n20111, n20112, n20113,
         n20114, n20115, n20116, n20117, n20118, n20119, n20120, n20121,
         n20122, n20123, n20124, n20125, n20126, n20127, n20128, n20129,
         n20130, n20131, n20132, n20133, n20134, n20135, n20136, n20137,
         n20138, n20139, n20140, n20141, n20142, n20143, n20144, n20145,
         n20146, n20147, n20148, n20149, n20150, n20151, n20152, n20153,
         n20154, n20155, n20156, n20157, n20158, n20159, n20160, n20161,
         n20162, n20163, n20164, n20165, n20166, n20167, n20168, n20169,
         n20170, n20171, n20172, n20173, n20174, n20175, n20176, n20177,
         n20178, n20179, n20180, n20181, n20182, n20183, n20184, n20185,
         n20186, n20187, n20188, n20189, n20190, n20191, n20192, n20193,
         n20194, n20195, n20196, n20197, n20198, n20199, n20200, n20201,
         n20202, n20203, n20204, n20205, n20206, n20207, n20208, n20209,
         n20210, n20211, n20212, n20213, n20214, n20215, n20216, n20217,
         n20218, n20219, n20220, n20221, n20222, n20223, n20224, n20225,
         n20226, n20227, n20228, n20229, n20230, n20231, n20232, n20233,
         n20234, n20235, n20236, n20237, n20238, n20239, n20240, n20241,
         n20242, n20243, n20244, n20245, n20246, n20247, n20248, n20249,
         n20250, n20251, n20252, n20253, n20254, n20255, n20256, n20257,
         n20258, n20259, n20260, n20261, n20262, n20263, n20264, n20265,
         n20266, n20267, n20268, n20269, n20270, n20271, n20272, n20273,
         n20274, n20275, n20276, n20277, n20278, n20279, n20280, n20281,
         n20282, n20283, n20284, n20285, n20286, n20287, n20288, n20289,
         n20290, n20291, n20292, n20293, n20294, n20295, n20296, n20297,
         n20298, n20299, n20300, n20301, n20302, n20303, n20304, n20305,
         n20306, n20307, n20308, n20309, n20310, n20311, n20312, n20313,
         n20314, n20315, n20316, n20317, n20318, n20319, n20320, n20321,
         n20322, n20323, n20324, n20325, n20326, n20327, n20328, n20329,
         n20330, n20331, n20332, n20333, n20334, n20335, n20336, n20337,
         n20338, n20339, n20340, n20341, n20342, n20343, n20344, n20345,
         n20346, n20347, n20348, n20349, n20350, n20351, n20352, n20353,
         n20354, n20355, n20356, n20357, n20358, n20359, n20360, n20361,
         n20362, n20363, n20364, n20365, n20366, n20367, n20368, n20369,
         n20370, n20371, n20372, n20373, n20374, n20375, n20376, n20377,
         n20378, n20379, n20380, n20381, n20382, n20383, n20384, n20385,
         n20386, n20387, n20388, n20389, n20390, n20391, n20392, n20393,
         n20394, n20395, n20396, n20397, n20398, n20399, n20400, n20401,
         n20402, n20403, n20404, n20405, n20406, n20407, n20408, n20409,
         n20410, n20411, n20412, n20413, n20414, n20415, n20416, n20417,
         n20418, n20419, n20420, n20421, n20422, n20423, n20424, n20425,
         n20426, n20427, n20428, n20429, n20430, n20431, n20432, n20433,
         n20434, n20435, n20436, n20437, n20438, n20439, n20440, n20441,
         n20442, n20443, n20444, n20445, n20446, n20447, n20448, n20449,
         n20450, n20451, n20452, n20453, n20454, n20455, n20456, n20457,
         n20458, n20459, n20460, n20461, n20462, n20463, n20464, n20465,
         n20466, n20467, n20468, n20469, n20470, n20471, n20472, n20473,
         n20474, n20475, n20476, n20477, n20478, n20479, n20480, n20481,
         n20482, n20483, n20484, n20485, n20486, n20487, n20488, n20489,
         n20490, n20491, n20492, n20493, n20494, n20495, n20496, n20497,
         n20498, n20499, n20500, n20501, n20502, n20503, n20504, n20505,
         n20506, n20507, n20508, n20509, n20510, n20511, n20512, n20513,
         n20514, n20515, n20516, n20517, n20518, n20519, n20520, n20521,
         n20522, n20523, n20524, n20525, n20526, n20527, n20528, n20529,
         n20530, n20531, n20532, n20533, n20534, n20535, n20536, n20537,
         n20538, n20539, n20540, n20541, n20542, n20543, n20544, n20545,
         n20546, n20547, n20548, n20549, n20550, n20551, n20552, n20553,
         n20554, n20555, n20556, n20557, n20558, n20559, n20560, n20561,
         n20562, n20563, n20564, n20565, n20566, n20567, n20568, n20569,
         n20570, n20571, n20572, n20573, n20574, n20575, n20576, n20577,
         n20578, n20579, n20580, n20581, n20582, n20583, n20584, n20585,
         n20586, n20587, n20588, n20589, n20590, n20591, n20592, n20593,
         n20594, n20595, n20596, n20597, n20598, n20599, n20600, n20601,
         n20602, n20603, n20604, n20605, n20606, n20607, n20608, n20609,
         n20610, n20611, n20612, n20613, n20614, n20615, n20616, n20617,
         n20618, n20619, n20620, n20621, n20622, n20623, n20624, n20625,
         n20626, n20627, n20628, n20629, n20630, n20631, n20632, n20633,
         n20634, n20635, n20636, n20637, n20638, n20639, n20640, n20641,
         n20642, n20643, n20644, n20645, n20646, n20647, n20648, n20649,
         n20650, n20651, n20652, n20653, n20654, n20655, n20656, n20657,
         n20658, n20659, n20660, n20661, n20662, n20663, n20664, n20665,
         n20666, n20667, n20668, n20669, n20670, n20671, n20672, n20673,
         n20674, n20675, n20676, n20677, n20678, n20679, n20680, n20681,
         n20682, n20683, n20684, n20685, n20686, n20687, n20688, n20689,
         n20690, n20691, n20692, n20693, n20694, n20695, n20696, n20697,
         n20698, n20699, n20700, n20701, n20702, n20703, n20704, n20705,
         n20706, n20707, n20708, n20709, n20710, n20711, n20712, n20713,
         n20714, n20715, n20716, n20717, n20718, n20719, n20720, n20721,
         n20722, n20723, n20724, n20725, n20726, n20727, n20728, n20729,
         n20730, n20731, n20732, n20733, n20734, n20735, n20736, n20737,
         n20738, n20739, n20740, n20741, n20742, n20743, n20744, n20745,
         n20746, n20747, n20748, n20749, n20750, n20751;

  dfrbp_1 _____________9_____436169 ( .D(n10140), .CLK(n10646), .RESET_B(reset), .Q(n20749), .Q_N(n10629) );
  dfrtp_1 ______________0_____ ( .D(n10592), .CLK(n10658), .RESET_B(reset), 
        .Q(n23668) );
  dfrtp_1 ________________ ( .D(n10591), .CLK(n10654), .RESET_B(reset), .Q(
        outData[31]) );
  dfrtp_1 _________________9_ ( .D(n10143), .CLK(n10659), .RESET_B(reset), .Q(
        n23934) );
  dfrtp_1 _____________9___0_ ( .D(n10589), .CLK(n10654), .RESET_B(reset), .Q(
        n23898) );
  dfrtp_1 ______________0___0_ ( .D(n10588), .CLK(n10655), .RESET_B(reset), 
        .Q(n12587) );
  dfrtp_1 ______________0_447459 ( .D(n10356), .CLK(n10669), .RESET_B(reset), 
        .Q(outData[30]) );
  dfrtp_1 ___________________436225 ( .D(n10142), .CLK(n10668), .RESET_B(reset), .Q(n23935) );
  dfrtp_1 _____________9___9_ ( .D(n10141), .CLK(n10659), .RESET_B(reset), .Q(
        n12318) );
  dfrtp_1 ______________0___9_ ( .D(n10510), .CLK(n10659), .RESET_B(reset), 
        .Q(_____90__34411) );
  dfrtp_1 ______________9_ ( .D(n10509), .CLK(n10659), .RESET_B(reset), .Q(
        outData[29]) );
  dfrtp_1 ___________________437994 ( .D(n10582), .CLK(n10664), .RESET_B(reset), .Q(n23773) );
  dfrtp_1 ___________________437479 ( .D(n10581), .CLK(n10665), .RESET_B(reset), .Q(n23786) );
  dfrtp_1 __________________438929 ( .D(n10580), .CLK(n10650), .RESET_B(reset), 
        .Q(n12487) );
  dfrbp_1 ___________________436660 ( .D(n10503), .CLK(n10647), .RESET_B(reset), .Q_N(n818) );
  dfrtp_1 ___________________436724 ( .D(n10419), .CLK(n10659), .RESET_B(reset), .Q(n12476) );
  dfrtp_1 _____________________0_443577 ( .D(n209), .CLK(n10659), .RESET_B(
        reset), .Q(n23995) );
  dfrtp_1 ___________________436233 ( .D(n10501), .CLK(n10668), .RESET_B(reset), .Q(n23997) );
  dfrtp_1 _____________9_____436188 ( .D(n10144), .CLK(n10651), .RESET_B(reset), .Q(n12467) );
  dfrtp_1 ______________0_____436018 ( .D(n10508), .CLK(n10659), .RESET_B(
        reset), .Q(__________0_______18822) );
  dfrbp_1 ________________436012 ( .D(n10507), .CLK(n10649), .RESET_B(reset), 
        .Q(outData[28]), .Q_N(n10612) );
  dfrtp_1 ___________________436299 ( .D(n10534), .CLK(n10668), .RESET_B(reset), .Q(n23936) );
  dfrbp_1 _____________9_____436193 ( .D(n10533), .CLK(n10646), .RESET_B(reset), .Q_N(n779) );
  dfrtp_1 _____________9_____436240 ( .D(n10303), .CLK(n10661), .RESET_B(reset), .Q(n12429) );
  dfrbp_1 _____________9_____436227 ( .D(n10511), .CLK(n10646), .RESET_B(reset), .Q_N(n811) );
  dfrtp_1 ______________0_____436025 ( .D(n10532), .CLK(n10668), .RESET_B(
        reset), .Q(______0__34499) );
  dfrtp_1 ________________436019 ( .D(n10531), .CLK(n10659), .RESET_B(reset), 
        .Q(n12412) );
  dfrtp_1 ___________________436292 ( .D(n10514), .CLK(n10667), .RESET_B(reset), .Q(n23937) );
  dfrtp_1 ___________________436357 ( .D(n10513), .CLK(n10667), .RESET_B(reset), .Q(n70) );
  dfrtp_1 ___________________436442 ( .D(n10512), .CLK(n10659), .RESET_B(reset), .Q(n69) );
  dfrtp_1 _____________9_____436201 ( .D(n10430), .CLK(n10659), .RESET_B(reset), .Q(n12580) );
  dfrtp_1 _____________9_____436314 ( .D(n10217), .CLK(n10659), .RESET_B(reset), .Q(n68) );
  dfrtp_1 _____________9_____436351 ( .D(n10544), .CLK(n10663), .RESET_B(reset), .Q(n23920) );
  dfrtp_1 ______________0_____436032 ( .D(n10427), .CLK(n10649), .RESET_B(
        reset), .Q(n23667) );
  dfrtp_1 ________________436024 ( .D(n10426), .CLK(n10650), .RESET_B(reset), 
        .Q(outData[26]) );
  dfrtp_1 ______________0_____436055 ( .D(n10543), .CLK(n10663), .RESET_B(
        reset), .Q(__________0_______18820) );
  dfrtp_1 ________________436040 ( .D(n10542), .CLK(n10663), .RESET_B(reset), 
        .Q(outData[24]) );
  dfrtp_1 ________________436049 ( .D(n10428), .CLK(n10659), .RESET_B(reset), 
        .Q(n12391) );
  dfrtp_1 ___________________436468 ( .D(n10545), .CLK(n10652), .RESET_B(reset), .Q(n756) );
  dfrtp_1 _________________0_436521 ( .D(n10469), .CLK(n10652), .RESET_B(reset), .Q(n12371) );
  dfrtp_1 ___________________436661 ( .D(n10539), .CLK(n10660), .RESET_B(reset), .Q(n23704) );
  dfrbp_1 _____________9_____436376 ( .D(n10538), .CLK(n10646), .RESET_B(reset), .Q_N(n771) );
  dfrtp_1 _____________9_____436510 ( .D(n10305), .CLK(n10652), .RESET_B(reset), .Q(n67) );
  dfrtp_1 _____________9_____436566 ( .D(n10304), .CLK(n10656), .RESET_B(reset), .Q(n12484) );
  dfrtp_1 ______________0_____436148 ( .D(n10537), .CLK(n10652), .RESET_B(
        reset), .Q(_____9___34413) );
  dfrtp_1 ________________436125 ( .D(n10536), .CLK(n10652), .RESET_B(reset), 
        .Q(outData[21]) );
  dfrtp_1 ______________0_____436107 ( .D(n10425), .CLK(n10659), .RESET_B(
        reset), .Q(__________0_______18818) );
  dfrtp_1 ________________436083 ( .D(n10424), .CLK(n10659), .RESET_B(reset), 
        .Q(n12426) );
  dfrtp_1 _________________9_438258 ( .D(n10196), .CLK(n10665), .RESET_B(reset), .Q(n23778) );
  dfrtp_1 ___________________437284 ( .D(n10598), .CLK(n10667), .RESET_B(reset), .Q(n66) );
  dfrtp_1 ___________________436682 ( .D(n10597), .CLK(n10667), .RESET_B(reset), .Q(n23885) );
  dfrtp_1 _________________9_436712 ( .D(n10596), .CLK(n10658), .RESET_B(reset), .Q(n12452) );
  dfrtp_1 ________________0_ ( .D(n10529), .CLK(n10667), .RESET_B(reset), .Q(
        n23882) );
  dfrbp_1 __________________ ( .D(n10553), .CLK(n10649), .RESET_B(reset), .Q(
        n10638), .Q_N(n698) );
  dfrtp_1 _____________9__9_ ( .D(n10574), .CLK(n10651), .RESET_B(reset), .Q(
        n12376) );
  dfrtp_1 ______________0___9_436203 ( .D(n10203), .CLK(n10660), .RESET_B(
        reset), .Q(n65) );
  dfrtp_1 ______________9_436179 ( .D(n10202), .CLK(n10661), .RESET_B(reset), 
        .Q(outData[19]) );
  dfrbp_1 _________________9_436572 ( .D(n10540), .CLK(n10649), .RESET_B(reset), .Q(n10633), .Q_N(n769) );
  dfrtp_1 _____________9___0_436272 ( .D(n10216), .CLK(n10663), .RESET_B(reset), .Q(n64) );
  dfrtp_1 ______________0___0_436144 ( .D(n10178), .CLK(n10661), .RESET_B(
        reset), .Q(__________0___0___18817) );
  dfrtp_1 ______________0_ ( .D(n10535), .CLK(n10661), .RESET_B(reset), .Q(
        outData[20]) );
  dfrtp_1 ______________0_____436437 ( .D(n10573), .CLK(n10656), .RESET_B(
        reset), .Q(______9__34498) );
  dfrtp_1 ________________436392 ( .D(n10572), .CLK(n10656), .RESET_B(reset), 
        .Q(n12413) );
  dfrtp_1 ___________________436861 ( .D(n10561), .CLK(n10656), .RESET_B(reset), .Q(n23943) );
  dfrtp_1 _____________9_____436654 ( .D(n10560), .CLK(n10655), .RESET_B(reset), .Q(n63) );
  dfrtp_1 _____________9_____436560 ( .D(n10307), .CLK(n10655), .RESET_B(reset), .Q(n12373) );
  dfrtp_1 _____________9_____436800 ( .D(n10556), .CLK(n10655), .RESET_B(reset), .Q(n62) );
  dfrtp_1 ______________0_____436284 ( .D(n10472), .CLK(n10655), .RESET_B(
        reset), .Q(n61) );
  dfrtp_1 ________________436253 ( .D(n10471), .CLK(n10655), .RESET_B(reset), 
        .Q(n12310) );
  dfrtp_1 ___________________436897 ( .D(n10504), .CLK(n10667), .RESET_B(reset), .Q(n60) );
  dfrtp_1 ___________________436903 ( .D(n10517), .CLK(n10659), .RESET_B(reset), .Q(n23803) );
  dfrtp_1 ___________________437047 ( .D(n10516), .CLK(n10667), .RESET_B(reset), .Q(n59) );
  dfrtp_1 ___________________436785 ( .D(n10515), .CLK(n10667), .RESET_B(reset), .Q(n23884) );
  dfrtp_1 ___________________436601 ( .D(n10211), .CLK(n10667), .RESET_B(reset), .Q(n12445) );
  dfrtp_1 ________________0_436608 ( .D(n10210), .CLK(n10657), .RESET_B(reset), 
        .Q(n12521) );
  dfrbp_1 _____________9__0_ ( .D(n10500), .CLK(n10647), .RESET_B(reset), .Q(
        n10639), .Q_N(n821) );
  dfrtp_1 _____________9____ ( .D(n10445), .CLK(n10657), .RESET_B(reset), .Q(
        n58) );
  dfrtp_1 ______________0_____436462 ( .D(n10555), .CLK(n10655), .RESET_B(
        reset), .Q(__________0_____) );
  dfrbp_1 ________________436428 ( .D(n10554), .CLK(n10647), .RESET_B(reset), 
        .Q(outData[12]), .Q_N(n10617) );
  dfrtp_1 ______________0_____436288 ( .D(n10559), .CLK(n10656), .RESET_B(
        reset), .Q(n57) );
  dfrtp_1 ________________436268 ( .D(n10558), .CLK(n10656), .RESET_B(reset), 
        .Q(outData[15]) );
  dfrtp_1 ___________________436809 ( .D(n10568), .CLK(n10666), .RESET_B(reset), .Q(n23945) );
  dfrtp_1 _________________0_436995 ( .D(n10570), .CLK(n10651), .RESET_B(reset), .Q(n23946) );
  dfrtp_1 _____________9_____436769 ( .D(n10308), .CLK(n10666), .RESET_B(reset), .Q(n23932) );
  dfrtp_1 ______________0_____436487 ( .D(n10478), .CLK(n10652), .RESET_B(
        reset), .Q(n56) );
  dfrbp_1 ________________436453 ( .D(n10477), .CLK(n10649), .RESET_B(reset), 
        .Q(outData[11]), .Q_N(n10611) );
  dfrtp_1 ______________0_____436326 ( .D(n10205), .CLK(n10667), .RESET_B(
        reset), .Q(n23666) );
  dfrtp_1 ________________436295 ( .D(n10571), .CLK(n10652), .RESET_B(reset), 
        .Q(outData[14]) );
  dfrtp_1 __________________437833 ( .D(n10520), .CLK(n10658), .RESET_B(reset), 
        .Q(n55) );
  dfrbp_1 ___________________437679 ( .D(n10462), .CLK(n10647), .RESET_B(reset), .Q(n23788), .Q_N(n10641) );
  dfrtp_1 _________________0_437788 ( .D(n10461), .CLK(n10646), .RESET_B(reset), .Q(n23789) );
  dfrtp_1 __________________437741 ( .D(n10460), .CLK(n10663), .RESET_B(reset), 
        .Q(n23856) );
  dfrtp_1 _________________0_437593 ( .D(n10458), .CLK(n10664), .RESET_B(reset), .Q(n23814) );
  dfrtp_1 __________________437648 ( .D(n10457), .CLK(n10664), .RESET_B(reset), 
        .Q(n23715) );
  dfrtp_1 __________________437482 ( .D(n10454), .CLK(n10658), .RESET_B(reset), 
        .Q(n23865) );
  dfrtp_1 __________________437425 ( .D(n10453), .CLK(n10650), .RESET_B(reset), 
        .Q(n23867) );
  dfrtp_1 _________________0_437325 ( .D(n10456), .CLK(n10658), .RESET_B(reset), .Q(n23857) );
  dfrtp_1 ________________9_437519 ( .D(n10455), .CLK(n10658), .RESET_B(reset), 
        .Q(n23767) );
  dfrtp_1 ________________9_ ( .D(n10575), .CLK(n10656), .RESET_B(reset), .Q(
        n12473) );
  dfrtp_1 _____________9___0_436659 ( .D(n10475), .CLK(n10651), .RESET_B(reset), .Q(n23928) );
  dfrtp_1 ______________0___0_436562 ( .D(n10474), .CLK(n10651), .RESET_B(
        reset), .Q(n23671) );
  dfrtp_1 ______________0_436494 ( .D(n10473), .CLK(n10651), .RESET_B(reset), 
        .Q(n12402) );
  dfrtp_1 __________________437202 ( .D(n10552), .CLK(n10658), .RESET_B(reset), 
        .Q(n54) );
  dfrtp_1 _____________9____437083 ( .D(n10481), .CLK(n10651), .RESET_B(reset), 
        .Q(n53) );
  dfrtp_1 ______________0__9_ ( .D(n10480), .CLK(n10651), .RESET_B(reset), .Q(
        n23672) );
  dfrtp_1 _____________9_ ( .D(n10479), .CLK(n10651), .RESET_B(reset), .Q(
        n12414) );
  dfrbp_1 __________________437600 ( .D(n10459), .CLK(n10648), .RESET_B(reset), 
        .Q(n23859), .Q_N(n10628) );
  dfrtp_1 __________________437556 ( .D(n10577), .CLK(n10666), .RESET_B(reset), 
        .Q(n23864) );
  dfrbp_1 __________________438414 ( .D(n10576), .CLK(n10646), .RESET_B(reset), 
        .Q(n20748) );
  dfrtp_1 __________________437163 ( .D(n10476), .CLK(n10651), .RESET_B(reset), 
        .Q(n52) );
  dfrbp_1 _____________9____436890 ( .D(n10451), .CLK(n10648), .RESET_B(reset), 
        .Q(n20750), .Q_N(n10631) );
  dfrtp_1 ______________0____ ( .D(n10442), .CLK(n10651), .RESET_B(reset), .Q(
        n51) );
  dfrtp_1 _______________ ( .D(n10441), .CLK(n10651), .RESET_B(reset), .Q(
        n12330) );
  dfrtp_1 __________________436986 ( .D(n10452), .CLK(n10656), .RESET_B(reset), 
        .Q(n23969) );
  dfrtp_1 _____________9____440211 ( .D(n10551), .CLK(n10656), .RESET_B(reset), 
        .Q(n12520) );
  dfrtp_1 ______________0____436697 ( .D(n10550), .CLK(n10650), .RESET_B(reset), .Q(n23669) );
  dfrtp_1 _______________436636 ( .D(n10549), .CLK(n10650), .RESET_B(reset), 
        .Q(outData[7]) );
  dfrtp_1 __________________437286 ( .D(n10528), .CLK(n10649), .RESET_B(reset), 
        .Q(n23924) );
  dfrtp_1 __________________438299 ( .D(n10152), .CLK(n10651), .RESET_B(reset), 
        .Q(n23925) );
  dfrtp_1 _____________9____440384 ( .D(n10527), .CLK(n10651), .RESET_B(reset), 
        .Q(n12547) );
  dfrtp_1 _____________9____440545 ( .D(n10209), .CLK(n10650), .RESET_B(reset), 
        .Q(n12549) );
  dfrtp_1 ______________0____439699 ( .D(n10526), .CLK(n10656), .RESET_B(reset), .Q(_____9___34419) );
  dfrbp_1 _______________439613 ( .D(n10525), .CLK(n10648), .RESET_B(reset), 
        .Q(outData[6]), .Q_N(n10619) );
  dfrtp_1 ______________0____439947 ( .D(n10448), .CLK(n10650), .RESET_B(reset), .Q(n50) );
  dfrbp_1 _______________439885 ( .D(n10447), .CLK(n10648), .RESET_B(reset), 
        .Q(n10604), .Q_N(outData[4]) );
  dfrtp_1 __________________439884 ( .D(n10524), .CLK(n10650), .RESET_B(reset), 
        .Q(n23706) );
  dfrtp_1 _____________9____440530 ( .D(n10208), .CLK(n10650), .RESET_B(reset), 
        .Q(n49) );
  dfrtp_1 ______________0____440093 ( .D(n10207), .CLK(n10651), .RESET_B(reset), .Q(n48) );
  dfrtp_1 _______________440017 ( .D(n10206), .CLK(n10650), .RESET_B(reset), 
        .Q(n12354) );
  dfrtp_1 ______________0____439790 ( .D(n10522), .CLK(n10650), .RESET_B(reset), .Q(n47) );
  dfrtp_1 _______________439722 ( .D(n10521), .CLK(n10650), .RESET_B(reset), 
        .Q(n12440) );
  dfrtp_1 __________________440748 ( .D(n10446), .CLK(n10656), .RESET_B(reset), 
        .Q(n23971) );
  dfrtp_1 _____________9____440715 ( .D(n10523), .CLK(n10657), .RESET_B(reset), 
        .Q(n46) );
  dfrtp_1 ______________0____440299 ( .D(n10177), .CLK(n10657), .RESET_B(reset), .Q(n45) );
  dfrtp_1 _______________440213 ( .D(n10176), .CLK(n10657), .RESET_B(reset), 
        .Q(n12308) );
  dfrtp_1 ______________0____441261 ( .D(n10444), .CLK(n10657), .RESET_B(reset), .Q(n44) );
  dfrtp_1 _______________441184 ( .D(n10443), .CLK(n10657), .RESET_B(reset), 
        .Q(n12506) );
  dfrtp_1 ______________0__0_ ( .D(n10499), .CLK(n10657), .RESET_B(reset), .Q(
        n12564) );
  dfrtp_1 ____0________________0_441664 ( .D(n10498), .CLK(n10657), .RESET_B(
        reset), .Q(n12384) );
  dfrtp_1 ____0_________________0_441885 ( .D(n10494), .CLK(n10657), .RESET_B(
        reset), .Q(n24035) );
  dfrbp_1 ____0__________________440749 ( .D(n10488), .CLK(n10649), .RESET_B(
        reset), .Q(n24029), .Q_N(n10610) );
  dfrtp_1 ____0__________________441339 ( .D(n10497), .CLK(n10657), .RESET_B(
        reset), .Q(n24032) );
  dfrtp_1 ____0__________________441547 ( .D(n10495), .CLK(n10657), .RESET_B(
        reset), .Q(n24026) );
  dfrtp_1 ____0___________________442326 ( .D(n10491), .CLK(n10657), .RESET_B(
        reset), .Q(n24023) );
  dfrtp_1 ____0__________________441828 ( .D(n10496), .CLK(n10657), .RESET_B(
        reset), .Q(n24024) );
  dfrtp_1 ____0__________________442437 ( .D(n10493), .CLK(n10658), .RESET_B(
        reset), .Q(n24030) );
  dfrtp_1 ____0__________________441591 ( .D(n10490), .CLK(n10658), .RESET_B(
        reset), .Q(n24028) );
  dfrtp_1 ____0________________9_ ( .D(n10492), .CLK(n10657), .RESET_B(reset), 
        .Q(n24025) );
  dfrtp_1 ____0__________________442180 ( .D(n10487), .CLK(n10658), .RESET_B(
        reset), .Q(n24033) );
  dfrtp_1 ____0__________________441604 ( .D(n10489), .CLK(n10657), .RESET_B(
        reset), .Q(n24027) );
  dfrtp_1 ____0___________________441638 ( .D(n10486), .CLK(n10658), .RESET_B(
        reset), .Q(n24031) );
  dfrbp_1 _______________________442355 ( .D(n10413), .CLK(n10647), .RESET_B(
        reset), .Q(n23982), .Q_N(n10622) );
  dfrtp_1 _______________________442613 ( .D(n10414), .CLK(n10660), .RESET_B(
        reset), .Q(n24003) );
  dfrtp_1 _______________________443184 ( .D(n10410), .CLK(n10660), .RESET_B(
        reset), .Q(n23983) );
  dfrtp_1 _____________________9_ ( .D(n10418), .CLK(n10660), .RESET_B(reset), 
        .Q(n24021) );
  dfrtp_1 _______________________440975 ( .D(n10412), .CLK(n10660), .RESET_B(
        reset), .Q(n24020) );
  dfrtp_1 _______________________441521 ( .D(n10417), .CLK(n10660), .RESET_B(
        reset), .Q(n23979) );
  dfrtp_1 _______________________442516 ( .D(n10415), .CLK(n10660), .RESET_B(
        reset), .Q(n24002) );
  dfrtp_1 _______________________442820 ( .D(n10411), .CLK(n10660), .RESET_B(
        reset), .Q(n24013) );
  dfrtp_1 _______________________442665 ( .D(n10416), .CLK(n10660), .RESET_B(
        reset), .Q(n24012) );
  dfrbp_1 _________________0_437850 ( .D(n10600), .CLK(n10649), .RESET_B(reset), .Q(n20745), .Q_N(n10635) );
  dfrtp_1 __________________437824 ( .D(n10601), .CLK(n10654), .RESET_B(reset), 
        .Q(n23840) );
  dfrtp_1 _________________9_437861 ( .D(n10223), .CLK(n10662), .RESET_B(reset), .Q(n23750) );
  dfrtp_1 _________________9_437953 ( .D(n10284), .CLK(n10662), .RESET_B(reset), .Q(n23765) );
  dfrtp_1 ___________________437882 ( .D(n10283), .CLK(n10653), .RESET_B(reset), .Q(n23736) );
  dfrtp_1 ___________________438034 ( .D(n10222), .CLK(n10653), .RESET_B(reset), .Q(n12351) );
  dfrtp_1 ___________________437952 ( .D(n10289), .CLK(n10653), .RESET_B(reset), .Q(n23694) );
  dfrtp_1 ___________________438000 ( .D(n10282), .CLK(n10653), .RESET_B(reset), .Q(n23875) );
  dfrtp_1 ___________________437898 ( .D(n10281), .CLK(n10662), .RESET_B(reset), .Q(n43) );
  dfrtp_1 ________________0_442232 ( .D(n10280), .CLK(n10662), .RESET_B(reset), 
        .Q(n42) );
  dfrtp_1 __________________441325 ( .D(n10584), .CLK(n10650), .RESET_B(reset), 
        .Q(n23877) );
  dfrtp_1 __________________437933 ( .D(n10226), .CLK(n10664), .RESET_B(reset), 
        .Q(n12518) );
  dfrbp_1 __________________437866 ( .D(n10227), .CLK(n10646), .RESET_B(reset), 
        .Q(n20747), .Q_N(n10630) );
  dfrtp_1 __________________441394 ( .D(n10583), .CLK(n10654), .RESET_B(reset), 
        .Q(n41) );
  dfrtp_1 __________________437837 ( .D(n10440), .CLK(n10664), .RESET_B(reset), 
        .Q(n23712) );
  dfrbp_1 __________________438684 ( .D(n10439), .CLK(n10649), .RESET_B(reset), 
        .Q(n23860), .Q_N(n10627) );
  dfrtp_1 _____________________0_443836 ( .D(n10438), .CLK(n10654), .RESET_B(
        reset), .Q(n24045) );
  dfrtp_1 _______________________442741 ( .D(n10378), .CLK(n10668), .RESET_B(
        reset), .Q(n24017) );
  dfrtp_1 ___________________437982 ( .D(n10286), .CLK(n10662), .RESET_B(reset), .Q(n23737) );
  dfrbp_1 ___________________438075 ( .D(n10288), .CLK(n10649), .RESET_B(reset), .Q(n23762), .Q_N(n10620) );
  dfrbp_1 ___________________444494 ( .D(n10285), .CLK(n10648), .RESET_B(reset), .Q(n20740), .Q_N(n10637) );
  dfrtp_1 ___________________438021 ( .D(n10291), .CLK(n10662), .RESET_B(reset), .Q(n23738) );
  dfrtp_1 ___________________444374 ( .D(n10290), .CLK(n10662), .RESET_B(reset), .Q(n40) );
  dfrtp_1 ___________________438038 ( .D(n10302), .CLK(n10662), .RESET_B(reset), .Q(n12513) );
  dfrbp_1 ___________________444436 ( .D(n10301), .CLK(n10647), .RESET_B(reset), .Q(n20742) );
  dfrtp_1 ___________________438082 ( .D(n10300), .CLK(n10662), .RESET_B(reset), .Q(n23740) );
  dfrtp_1 ___________________438220 ( .D(n10299), .CLK(n10663), .RESET_B(reset), .Q(n23760) );
  dfrtp_1 ___________________438259 ( .D(n10298), .CLK(n10673), .RESET_B(reset), .Q(n23741) );
  dfrtp_1 ___________________438353 ( .D(n10219), .CLK(n10673), .RESET_B(reset), .Q(n12485) );
  dfrtp_1 _________________0_438260 ( .D(n10295), .CLK(n10673), .RESET_B(reset), .Q(n23727) );
  dfrtp_1 _____________________0_442818 ( .D(n10468), .CLK(n10652), .RESET_B(
        reset), .Q(n23903) );
  dfrtp_1 _____________________9_441409 ( .D(n10407), .CLK(n10652), .RESET_B(
        reset), .Q(n23992) );
  dfrtp_1 _______________________441590 ( .D(n10399), .CLK(n10653), .RESET_B(
        reset), .Q(n24000) );
  dfrtp_1 ______________________0_441637 ( .D(n10467), .CLK(n10652), .RESET_B(
        reset), .Q(n23991) );
  dfrtp_1 _______________________441300 ( .D(n10405), .CLK(n10652), .RESET_B(
        reset), .Q(n24008) );
  dfrtp_1 _______________________441488 ( .D(n10409), .CLK(n10652), .RESET_B(
        reset), .Q(n23972) );
  dfrbp_1 _______________________441946 ( .D(n10400), .CLK(n10648), .RESET_B(
        reset), .Q(n24009), .Q_N(n10626) );
  dfrbp_1 _______________________441257 ( .D(n10402), .CLK(n10649), .RESET_B(
        reset), .Q(n23998), .Q_N(n10621) );
  dfrbp_1 _______________________441062 ( .D(n10408), .CLK(n10648), .RESET_B(
        reset), .Q(n10624), .Q_N(n1678) );
  dfrtp_1 _______________________441485 ( .D(n10403), .CLK(n10652), .RESET_B(
        reset), .Q(n23999) );
  dfrbp_1 ________________________441694 ( .D(n10404), .CLK(n10649), .RESET_B(
        reset), .Q(n23990) );
  dfrtp_1 _______________________441679 ( .D(n10406), .CLK(n10652), .RESET_B(
        reset), .Q(n24001) );
  dfrtp_1 ________________________441542 ( .D(n10401), .CLK(n10653), .RESET_B(
        reset), .Q(n23970) );
  dfrtp_1 _____________________0_ ( .D(n10450), .CLK(n10658), .RESET_B(reset), 
        .Q(n12297) );
  dfrbp_1 ________________________442568 ( .D(n10398), .CLK(n10648), .RESET_B(
        reset), .Q(n23964), .Q_N(n10616) );
  dfrtp_1 _____________________9_442564 ( .D(n10395), .CLK(n10653), .RESET_B(
        reset), .Q(n23974) );
  dfrtp_1 ________________________443009 ( .D(n10449), .CLK(n10652), .RESET_B(
        reset), .Q(n23960) );
  dfrtp_1 ______________________0_ ( .D(n10393), .CLK(n10653), .RESET_B(reset), 
        .Q(n23962) );
  dfrtp_1 _______________________440974 ( .D(n10389), .CLK(n10653), .RESET_B(
        reset), .Q(n23978) );
  dfrtp_1 _______________________442664 ( .D(n10388), .CLK(n10653), .RESET_B(
        reset), .Q(n24005) );
  dfrbp_1 _______________________ ( .D(n215), .CLK(n10647), .RESET_B(reset), 
        .Q(n23977) );
  dfrtp_1 _______________________442478 ( .D(n10390), .CLK(n10653), .RESET_B(
        reset), .Q(n23975) );
  dfrtp_1 ________________________ ( .D(n10311), .CLK(n10653), .RESET_B(reset), 
        .Q(n23961) );
  dfrtp_1 _______________________442712 ( .D(n10397), .CLK(n10653), .RESET_B(
        reset), .Q(n24006) );
  dfrtp_1 _______________________442480 ( .D(n10392), .CLK(n10653), .RESET_B(
        reset), .Q(n23976) );
  dfrbp_1 _______________________442519 ( .D(n10391), .CLK(n10648), .RESET_B(
        reset), .Q(n24004), .Q_N(n10605) );
  dfrbp_1 _______________________442400 ( .D(n10394), .CLK(n10648), .RESET_B(
        reset), .Q(n24007), .Q_N(n10615) );
  dfrtp_1 _______________________442399 ( .D(n10387), .CLK(n10654), .RESET_B(
        reset), .Q(n24038) );
  dfrtp_1 _______________________441545 ( .D(n10379), .CLK(n10654), .RESET_B(
        reset), .Q(n23986) );
  dfrtp_1 _____________________9_442612 ( .D(n10385), .CLK(n10654), .RESET_B(
        reset), .Q(n12472) );
  dfrtp_1 _______________________442794 ( .D(n10381), .CLK(n10654), .RESET_B(
        reset), .Q(n24040) );
  dfrtp_1 _______________________443218 ( .D(n10383), .CLK(n10654), .RESET_B(
        reset), .Q(n24042) );
  dfrtp_1 ________________________441354 ( .D(n10384), .CLK(n10654), .RESET_B(
        reset), .Q(n12355) );
  dfrtp_1 ______________________0_441649 ( .D(n198), .CLK(n10654), .RESET_B(
        reset), .Q(n12316) );
  dfrbp_1 _______________________442710 ( .D(n10386), .CLK(n10646), .RESET_B(
        reset), .Q(n24039), .Q_N(n10636) );
  dfrtp_1 _______________________442517 ( .D(n10380), .CLK(n10671), .RESET_B(
        reset), .Q(n24047) );
  dfrtp_1 _______________________442566 ( .D(n10382), .CLK(n10654), .RESET_B(
        reset), .Q(n24046) );
  dfrtp_1 ________________________442115 ( .D(n10396), .CLK(n10653), .RESET_B(
        reset), .Q(n23963) );
  dfrtp_1 __________________440604 ( .D(n10309), .CLK(n10672), .RESET_B(reset), 
        .Q(n39) );
  dfrbp_1 __________________439906 ( .D(n10276), .CLK(n10648), .RESET_B(reset), 
        .Q_N(n2047) );
  dfrtp_1 __________________439405 ( .D(n10271), .CLK(n10668), .RESET_B(reset), 
        .Q(n23711) );
  dfrtp_1 __________________439795 ( .D(n10483), .CLK(n10668), .RESET_B(reset), 
        .Q(n23850) );
  dfrtp_1 _____________________0_439590 ( .D(n10482), .CLK(n10668), .RESET_B(
        reset), .Q(n23922) );
  dfrtp_1 ______________________0_442518 ( .D(n10369), .CLK(n10668), .RESET_B(
        reset), .Q(n23873) );
  dfrtp_1 _____________________9_441621 ( .D(n10374), .CLK(n10668), .RESET_B(
        reset), .Q(n23871) );
  dfrtp_1 _______________________441805 ( .D(n10370), .CLK(n10669), .RESET_B(
        reset), .Q(n24037) );
  dfrtp_1 _______________________442181 ( .D(n10368), .CLK(n10669), .RESET_B(
        reset), .Q(n23894) );
  dfrtp_1 _______________________442479 ( .D(n10367), .CLK(n10669), .RESET_B(
        reset), .Q(n23895) );
  dfrtp_1 _______________________441806 ( .D(n10371), .CLK(n10668), .RESET_B(
        reset), .Q(n23893) );
  dfrtp_1 _______________________441817 ( .D(n10365), .CLK(n10669), .RESET_B(
        reset), .Q(n23892) );
  dfrtp_1 ________________________441981 ( .D(n10373), .CLK(n10668), .RESET_B(
        reset), .Q(n23872) );
  dfrtp_1 _______________________442143 ( .D(n10366), .CLK(n10669), .RESET_B(
        reset), .Q(n23836) );
  dfrtp_1 ________________________442045 ( .D(n10364), .CLK(n10669), .RESET_B(
        reset), .Q(n24036) );
  dfrbp_1 _______________________442081 ( .D(n10372), .CLK(n10646), .RESET_B(
        reset), .Q(n23837), .Q_N(n10614) );
  dfrtp_1 _______________________442713 ( .D(n10363), .CLK(n10669), .RESET_B(
        reset), .Q(n23838) );
  dfrtp_1 ____0________________0_ ( .D(n10587), .CLK(n10655), .RESET_B(reset), 
        .Q(n12558) );
  dfrtp_1 ____0__________________442210 ( .D(n10362), .CLK(n10669), .RESET_B(
        reset), .Q(n24057) );
  dfrtp_1 ____0___________________ ( .D(n10357), .CLK(n10669), .RESET_B(reset), 
        .Q(n24052) );
  dfrbp_1 ____0__________________442268 ( .D(n10377), .CLK(n10647), .RESET_B(
        reset), .Q(n20751), .Q_N(n10618) );
  dfrtp_1 ____0___________________441031 ( .D(n10375), .CLK(n10655), .RESET_B(
        reset), .Q(n24051) );
  dfrtp_1 ____0__________________442569 ( .D(n10355), .CLK(n10669), .RESET_B(
        reset), .Q(n24061) );
  dfrtp_1 ____0__________________440670 ( .D(n10352), .CLK(n10670), .RESET_B(
        reset), .Q(n38) );
  dfrtp_1 ____0__________________441032 ( .D(n10359), .CLK(n10669), .RESET_B(
        reset), .Q(n24053) );
  dfrtp_1 ____0_________________0_ ( .D(n10361), .CLK(n10669), .RESET_B(reset), 
        .Q(n24048) );
  dfrbp_1 ____0__________________442663 ( .D(n10354), .CLK(n10647), .RESET_B(
        reset), .Q(n24056), .Q_N(n10613) );
  dfrtp_1 ____0________________9_442254 ( .D(n10353), .CLK(n10669), .RESET_B(
        reset), .Q(n24054) );
  dfrtp_1 ____0__________________ ( .D(n10358), .CLK(n10655), .RESET_B(reset), 
        .Q(n24059) );
  dfrtp_1 ____0___________________442354 ( .D(n10360), .CLK(n10669), .RESET_B(
        reset), .Q(n24062) );
  dfrtp_1 ____0__________________442356 ( .D(n10351), .CLK(n10670), .RESET_B(
        reset), .Q(n24058) );
  dfrtp_1 ____0___________________441126 ( .D(n10376), .CLK(n10655), .RESET_B(
        reset), .Q(n24055) );
  dfrtp_1 _____________0_ ( .D(n10350), .CLK(n10669), .RESET_B(reset), .Q(
        n12464) );
  dfrtp_1 ________________9_442357 ( .D(n10342), .CLK(n10670), .RESET_B(reset), 
        .Q(n23958) );
  dfrtp_1 __________________445195 ( .D(n10345), .CLK(n10670), .RESET_B(reset), 
        .Q(n12393) );
  dfrbp_1 __________________443904 ( .D(n10344), .CLK(n10647), .RESET_B(reset), 
        .Q(n10606), .Q_N(n1965) );
  dfrtp_1 __________________443074 ( .D(n10343), .CLK(n10670), .RESET_B(reset), 
        .Q(n12340) );
  dfrtp_1 __________________442913 ( .D(n10330), .CLK(n10671), .RESET_B(reset), 
        .Q(n23951) );
  dfrtp_1 __________________444880 ( .D(n10332), .CLK(n10671), .RESET_B(reset), 
        .Q(n12299) );
  dfrtp_1 __________________443811 ( .D(n10329), .CLK(n10671), .RESET_B(reset), 
        .Q(n23953) );
  dfrtp_1 _________________9_444058 ( .D(n10294), .CLK(n10673), .RESET_B(reset), .Q(n12479) );
  dfrtp_1 __________________443493 ( .D(n10331), .CLK(n10671), .RESET_B(reset), 
        .Q(n12320) );
  dfrtp_1 ___________________442912 ( .D(n10297), .CLK(n10673), .RESET_B(reset), .Q(n2029) );
  dfrtp_1 _________________0_447808 ( .D(n10296), .CLK(n10673), .RESET_B(reset), .Q(n23728) );
  dfrtp_1 __________________442883 ( .D(n10336), .CLK(n10671), .RESET_B(reset), 
        .Q(n23948) );
  dfrtp_1 __________________444879 ( .D(n10335), .CLK(n10672), .RESET_B(reset), 
        .Q(n12302) );
  dfrtp_1 __________________444159 ( .D(n10334), .CLK(n10672), .RESET_B(reset), 
        .Q(n12319) );
  dfrtp_1 ________________0_443182 ( .D(n10333), .CLK(n10672), .RESET_B(reset), 
        .Q(n23959) );
  dfrtp_1 __________________443260 ( .D(n10317), .CLK(n10670), .RESET_B(reset), 
        .Q(n12392) );
  dfrtp_1 __________________442742 ( .D(n10321), .CLK(n10670), .RESET_B(reset), 
        .Q(n23981) );
  dfrtp_1 __________________449255 ( .D(n10316), .CLK(n10670), .RESET_B(reset), 
        .Q(n37) );
  dfrtp_1 __________________444745 ( .D(n10320), .CLK(n10670), .RESET_B(reset), 
        .Q(n12394) );
  dfrtp_1 __________________444156 ( .D(n10319), .CLK(n10670), .RESET_B(reset), 
        .Q(n23828) );
  dfrtp_1 __________________443762 ( .D(n10318), .CLK(n10670), .RESET_B(reset), 
        .Q(n23987) );
  dfrtp_1 _______________0_ ( .D(n10347), .CLK(n10670), .RESET_B(reset), .Q(
        n24019) );
  dfrbp_1 _________________442770 ( .D(n10346), .CLK(n10647), .RESET_B(reset), 
        .Q(n24015), .Q_N(n10609) );
  dfrtp_1 _________________444216 ( .D(n10349), .CLK(n10670), .RESET_B(reset), 
        .Q(n12408) );
  dfrtp_1 _________________443620 ( .D(n10348), .CLK(n10670), .RESET_B(reset), 
        .Q(n12331) );
  dfrtp_1 _________________445093 ( .D(n10341), .CLK(n10671), .RESET_B(reset), 
        .Q(n12333) );
  dfrtp_1 _________________443665 ( .D(n10340), .CLK(n10671), .RESET_B(reset), 
        .Q(n23993) );
  dfrtp_1 __________________450844 ( .D(n10603), .CLK(n10672), .RESET_B(reset), 
        .Q(n23829) );
  dfrbp_1 _________________444743 ( .D(n10339), .CLK(n10648), .RESET_B(reset), 
        .Q(n24011), .Q_N(n10608) );
  dfrtp_1 ________________0_450796 ( .D(n10338), .CLK(n10671), .RESET_B(reset), 
        .Q(n36) );
  dfrtp_1 _________________444742 ( .D(n10337), .CLK(n10671), .RESET_B(reset), 
        .Q(n24022) );
  dfrtp_1 ________________0_440938 ( .D(n10279), .CLK(n10653), .RESET_B(reset), 
        .Q(n23876) );
  dfrtp_1 _________________ ( .D(n10324), .CLK(n10671), .RESET_B(reset), .Q(
        n12401) );
  dfrtp_1 __________________440868 ( .D(n10602), .CLK(n10672), .RESET_B(reset), 
        .Q(n23686) );
  dfrtp_1 __________________442795 ( .D(n10322), .CLK(n10671), .RESET_B(reset), 
        .Q(n23985) );
  dfrtp_1 ________________0_444744 ( .D(n10328), .CLK(n10671), .RESET_B(reset), 
        .Q(n12388) );
  dfrtp_1 __________________444157 ( .D(n10325), .CLK(n10671), .RESET_B(reset), 
        .Q(n35) );
  dfrtp_1 _______________9_ ( .D(n10327), .CLK(n10670), .RESET_B(reset), .Q(
        n12305) );
  dfrtp_1 __________________443528 ( .D(n10326), .CLK(n10671), .RESET_B(reset), 
        .Q(n34) );
  dfrtp_1 __________________439259 ( .D(n10230), .CLK(n10663), .RESET_B(reset), 
        .Q(n23853) );
  dfrtp_1 __________________438797 ( .D(n10160), .CLK(n10654), .RESET_B(reset), 
        .Q(n12510) );
  dfrtp_1 __________________450831 ( .D(n10323), .CLK(n10671), .RESET_B(reset), 
        .Q(n12586) );
  dfrtp_1 __________________440729 ( .D(n10310), .CLK(n10672), .RESET_B(reset), 
        .Q(n12584) );
  dfrtp_1 __________________440510 ( .D(n10485), .CLK(n10672), .RESET_B(reset), 
        .Q(n1144) );
  dfrtp_1 __________________440554 ( .D(n10278), .CLK(n10673), .RESET_B(reset), 
        .Q(n2045) );
  dfrtp_1 __________________440348 ( .D(n10233), .CLK(n10672), .RESET_B(reset), 
        .Q(n33) );
  dfrtp_1 __________________438441 ( .D(n10157), .CLK(n10654), .RESET_B(reset), 
        .Q(n23709) );
  dfrtp_1 __________________440224 ( .D(n10484), .CLK(n10673), .RESET_B(reset), 
        .Q(n32) );
  dfrtp_1 ________________0_443958 ( .D(n10315), .CLK(n10672), .RESET_B(reset), 
        .Q(n23949) );
  dfrbp_1 ________________9_447525 ( .D(n10314), .CLK(n10649), .RESET_B(reset), 
        .Q(n23950), .Q_N(n10607) );
  dfrtp_1 __________________446037 ( .D(n10313), .CLK(n10672), .RESET_B(reset), 
        .Q(n23938) );
  dfrtp_1 __________________445962 ( .D(n10312), .CLK(n10672), .RESET_B(reset), 
        .Q(n12380) );
  dfrtp_1 ___________________437924 ( .D(n10224), .CLK(n10662), .RESET_B(reset), .Q(n31) );
  dfrtp_1 ______________0_____436044 ( .D(n10145), .CLK(n10663), .RESET_B(
        reset), .Q(n23870) );
  dfrtp_1 ________________436033 ( .D(n10541), .CLK(n10663), .RESET_B(reset), 
        .Q(outData[25]) );
  dfrtp_1 ______________0_____436229 ( .D(n10204), .CLK(n10656), .RESET_B(
        reset), .Q(n30) );
  dfrtp_1 ______________0_____436244 ( .D(n10566), .CLK(n10655), .RESET_B(
        reset), .Q(n29) );
  dfrtp_1 ________________436207 ( .D(n10565), .CLK(n10655), .RESET_B(reset), 
        .Q(n12346) );
  dfrtp_1 ________________436202 ( .D(n10470), .CLK(n10656), .RESET_B(reset), 
        .Q(outData[18]) );
  dfrtp_1 __________________440422 ( .D(n10269), .CLK(n10673), .RESET_B(reset), 
        .Q(n12486) );
  dfrtp_1 __________________440172 ( .D(n10270), .CLK(n10672), .RESET_B(reset), 
        .Q(n12451) );
  dfrtp_1 __________________439636 ( .D(n10274), .CLK(n10658), .RESET_B(reset), 
        .Q(n28) );
  dfrtp_1 __________________446645 ( .D(n10273), .CLK(n10670), .RESET_B(reset), 
        .Q(n12450) );
  dfrbp_1 __________________439637 ( .D(n10275), .CLK(n10648), .RESET_B(reset), 
        .Q(n23833), .Q_N(n10645) );
  dfrtp_1 __________________439905 ( .D(n10466), .CLK(n10672), .RESET_B(reset), 
        .Q(n23831) );
  dfrtp_1 __________________439712 ( .D(n10465), .CLK(n10672), .RESET_B(reset), 
        .Q(n23845) );
  dfrtp_1 _________________0_439638 ( .D(n10266), .CLK(n10674), .RESET_B(reset), .Q(n27) );
  dfrtp_1 _________________0_439515 ( .D(n10268), .CLK(n10674), .RESET_B(reset), .Q(n26) );
  dfrtp_1 ________________9_439258 ( .D(n10267), .CLK(n10674), .RESET_B(reset), 
        .Q(n12583) );
  dfrtp_1 ________________9_439794 ( .D(n10238), .CLK(n10650), .RESET_B(reset), 
        .Q(n23830) );
  dfrtp_1 ________________9_439584 ( .D(n10237), .CLK(n10673), .RESET_B(reset), 
        .Q(n25) );
  dfrtp_1 _________________9_438507 ( .D(n10239), .CLK(n10673), .RESET_B(reset), .Q(n24) );
  dfrtp_1 ___________________438322 ( .D(n10244), .CLK(n10673), .RESET_B(reset), .Q(n23743) );
  dfrtp_1 _________________9_438338 ( .D(n10246), .CLK(n10673), .RESET_B(reset), .Q(n23742) );
  dfrbp_1 ___________________447225 ( .D(n10245), .CLK(n10647), .RESET_B(reset), .Q(n20741), .Q_N(n10642) );
  dfrtp_1 ___________________438542 ( .D(n10243), .CLK(n10673), .RESET_B(reset), .Q(n23758) );
  dfrtp_1 ___________________444215 ( .D(n10242), .CLK(n10673), .RESET_B(reset), .Q(n23730) );
  dfrtp_1 ___________________447193 ( .D(n10241), .CLK(n10673), .RESET_B(reset), .Q(n12516) );
  dfrbp_1 ___________________438701 ( .D(n10240), .CLK(n10647), .RESET_B(reset), .Q(n20743), .Q_N(n10640) );
  dfrtp_1 _________________0_438413 ( .D(n10220), .CLK(n10663), .RESET_B(reset), .Q(n23759) );
  dfrtp_1 ___________________438531 ( .D(n10262), .CLK(n10674), .RESET_B(reset), .Q(n23682) );
  dfrbp_1 ___________________438775 ( .D(n10261), .CLK(n10646), .RESET_B(reset), .Q_N(n2056) );
  dfrtp_1 ___________________443576 ( .D(n10260), .CLK(n10674), .RESET_B(reset), .Q(n12480) );
  dfrtp_1 ___________________438764 ( .D(n10258), .CLK(n10662), .RESET_B(reset), .Q(n23753) );
  dfrtp_1 ___________________438869 ( .D(n10259), .CLK(n10674), .RESET_B(reset), .Q(n23745) );
  dfrtp_1 ___________________447224 ( .D(n10257), .CLK(n10661), .RESET_B(reset), .Q(n12475) );
  dfrtp_1 ___________________438946 ( .D(n10256), .CLK(n10661), .RESET_B(reset), .Q(n23757) );
  dfrtp_1 ___________________439051 ( .D(n10255), .CLK(n10674), .RESET_B(reset), .Q(n23746) );
  dfrtp_1 ___________________439023 ( .D(n10254), .CLK(n10674), .RESET_B(reset), .Q(n23) );
  dfrtp_1 ___________________439222 ( .D(n10253), .CLK(n10674), .RESET_B(reset), .Q(n23747) );
  dfrtp_1 ___________________444158 ( .D(n10252), .CLK(n10674), .RESET_B(reset), .Q(n22) );
  dfrtp_1 ___________________447045 ( .D(n10247), .CLK(n10674), .RESET_B(reset), .Q(n23733) );
  dfrtp_1 ___________________439163 ( .D(n10248), .CLK(n10674), .RESET_B(reset), .Q(n23683) );
  dfrtp_1 ___________________439002 ( .D(n10251), .CLK(n10674), .RESET_B(reset), .Q(n23748) );
  dfrtp_1 ___________________443007 ( .D(n10250), .CLK(n10674), .RESET_B(reset), .Q(n12441) );
  dfrtp_1 ___________________439444 ( .D(n10265), .CLK(n10674), .RESET_B(reset), .Q(n12481) );
  dfrtp_1 ___________________439416 ( .D(n10264), .CLK(n10651), .RESET_B(reset), .Q(n23754) );
  dfrtp_1 _________________0_442709 ( .D(n10263), .CLK(n10674), .RESET_B(reset), .Q(n23725) );
  dfrtp_1 ___________________439330 ( .D(n10249), .CLK(n10664), .RESET_B(reset), .Q(n23756) );
  dfrtp_1 ___________________438622 ( .D(n10185), .CLK(n10662), .RESET_B(reset), .Q(n23780) );
  dfrtp_1 ___________________438683 ( .D(n10188), .CLK(n10660), .RESET_B(reset), .Q(n23781) );
  dfrtp_1 ___________________438754 ( .D(n10187), .CLK(n10661), .RESET_B(reset), .Q(n23696) );
  dfrtp_1 ___________________438848 ( .D(n10186), .CLK(n10661), .RESET_B(reset), .Q(n23691) );
  dfrtp_1 __________________440016 ( .D(n10272), .CLK(n10672), .RESET_B(reset), 
        .Q(n23843) );
  dfrtp_1 __________________440202 ( .D(n10235), .CLK(n10673), .RESET_B(reset), 
        .Q(n21) );
  dfrtp_1 __________________439614 ( .D(n10586), .CLK(n10663), .RESET_B(reset), 
        .Q(n12517) );
  dfrtp_1 __________________439105 ( .D(n10228), .CLK(n10663), .RESET_B(reset), 
        .Q(n23854) );
  dfrtp_1 __________________439781 ( .D(n10585), .CLK(n10663), .RESET_B(reset), 
        .Q(n23878) );
  dfrtp_1 ________________0_441544 ( .D(n10232), .CLK(n10662), .RESET_B(reset), 
        .Q(n20) );
  dfrtp_1 ________________0_441930 ( .D(n10225), .CLK(n10663), .RESET_B(reset), 
        .Q(n23880) );
  dfrtp_1 __________________440825 ( .D(n10159), .CLK(n10665), .RESET_B(reset), 
        .Q(n19) );
  dfrtp_1 __________________438604 ( .D(n10234), .CLK(n10656), .RESET_B(reset), 
        .Q(n23848) );
  dfrtp_1 ___________________438551 ( .D(n10463), .CLK(n10656), .RESET_B(reset), .Q(n23782) );
  dfrtp_1 _________________0_438977 ( .D(n10236), .CLK(n10672), .RESET_B(reset), .Q(n12430) );
  dfrtp_1 ________________9_438821 ( .D(n10464), .CLK(n10674), .RESET_B(reset), 
        .Q(n18) );
  dfrtp_1 ________________9_437762 ( .D(n10229), .CLK(n10658), .RESET_B(reset), 
        .Q(n23714) );
  dfrbp_1 __________________439688 ( .D(n10277), .CLK(n10647), .RESET_B(reset), 
        .Q_N(n2046) );
  dfrtp_1 __________________439423 ( .D(n10231), .CLK(n10651), .RESET_B(reset), 
        .Q(n2074) );
  dfrtp_1 __________________438813 ( .D(n10579), .CLK(n10650), .RESET_B(reset), 
        .Q(n23861) );
  dfrtp_1 ________________0_441264 ( .D(n10158), .CLK(n10650), .RESET_B(reset), 
        .Q(n23687) );
  dfrtp_1 __________________440374 ( .D(n10578), .CLK(n10666), .RESET_B(reset), 
        .Q(n23869) );
  dfrbp_1 ___________________438236 ( .D(n10195), .CLK(n10648), .RESET_B(reset), .Q(n23784), .Q_N(n10643) );
  dfrbp_1 ___________________438357 ( .D(n10194), .CLK(n10647), .RESET_B(reset), .Q(n23779), .Q_N(n10634) );
  dfrtp_1 ___________________438447 ( .D(n10197), .CLK(n10665), .RESET_B(reset), .Q(n23783) );
  dfrbp_1 ___________________438198 ( .D(n10221), .CLK(n10648), .RESET_B(reset), .Q(n20744) );
  dfrtp_1 ___________________437995 ( .D(n10200), .CLK(n10665), .RESET_B(reset), .Q(n23774) );
  dfrtp_1 ___________________438108 ( .D(n10199), .CLK(n10665), .RESET_B(reset), .Q(n23775) );
  dfrbp_1 ___________________438156 ( .D(n10198), .CLK(n10649), .RESET_B(reset), .Q(n20746), .Q_N(n10632) );
  dfrtp_1 _________________0_438214 ( .D(n10201), .CLK(n10665), .RESET_B(reset), .Q(n17) );
  dfrtp_1 ___________________437565 ( .D(n10189), .CLK(n10665), .RESET_B(reset), .Q(n23796) );
  dfrtp_1 _________________0_437485 ( .D(n10192), .CLK(n10665), .RESET_B(reset), .Q(n23795) );
  dfrtp_1 ___________________437394 ( .D(n10191), .CLK(n10665), .RESET_B(reset), .Q(n23787) );
  dfrbp_1 ___________________437500 ( .D(n10190), .CLK(n10646), .RESET_B(reset), .Q(n23766), .Q_N(n10625) );
  dfrtp_1 ___________________437102 ( .D(n10155), .CLK(n10650), .RESET_B(reset), .Q(n12372) );
  dfrtp_1 ___________________436725 ( .D(n10212), .CLK(n10667), .RESET_B(reset), .Q(n12446) );
  dfrtp_1 ___________________437109 ( .D(n10154), .CLK(n10666), .RESET_B(reset), .Q(n23815) );
  dfrbp_1 __________________438710 ( .D(n10153), .CLK(n10646), .RESET_B(reset), 
        .Q_N(n2122) );
  dfrtp_1 __________________438499 ( .D(n10156), .CLK(n10665), .RESET_B(reset), 
        .Q(n23863) );
  dfrtp_1 ___________________438090 ( .D(n10293), .CLK(n10662), .RESET_B(reset), .Q(n23693) );
  dfrtp_1 ___________________438103 ( .D(n10292), .CLK(n10662), .RESET_B(reset), .Q(n23763) );
  dfrtp_1 ___________________444616 ( .D(n10287), .CLK(n10662), .RESET_B(reset), .Q(n23720) );
  dfrtp_1 ___________________437927 ( .D(n10423), .CLK(n10663), .RESET_B(reset), .Q(n16) );
  dfrtp_1 ___________________437867 ( .D(n10422), .CLK(n10664), .RESET_B(reset), .Q(n23681) );
  dfrtp_1 ___________________437421 ( .D(n10421), .CLK(n10665), .RESET_B(reset), .Q(n23797) );
  dfrtp_1 ___________________437914 ( .D(n10506), .CLK(n10666), .RESET_B(reset), .Q(n23772) );
  dfrtp_1 ___________________437886 ( .D(n10150), .CLK(n10666), .RESET_B(reset), .Q(n15) );
  dfrtp_1 __________________437812 ( .D(n10519), .CLK(n10663), .RESET_B(reset), 
        .Q(n23851) );
  dfrtp_1 ___________________437304 ( .D(n10518), .CLK(n10666), .RESET_B(reset), .Q(n23799) );
  dfrtp_1 ___________________437393 ( .D(n10193), .CLK(n10666), .RESET_B(reset), .Q(n12579) );
  dfrtp_1 ___________________436969 ( .D(n10420), .CLK(n10667), .RESET_B(reset), .Q(n23804) );
  dfrtp_1 ___________________436743 ( .D(n10502), .CLK(n10668), .RESET_B(reset), .Q(n12522) );
  dfrtp_1 _________________9_437860 ( .D(n10149), .CLK(n10666), .RESET_B(reset), .Q(n23770) );
  dfrtp_1 _________________0_437798 ( .D(n10148), .CLK(n10666), .RESET_B(reset), .Q(n23680) );
  dfrtp_1 _________________0_437218 ( .D(n10147), .CLK(n10667), .RESET_B(reset), .Q(n23721) );
  dfrtp_1 _________________9_437326 ( .D(n10146), .CLK(n10667), .RESET_B(reset), .Q(n23769) );
  dfrtp_1 ___________________437362 ( .D(n10505), .CLK(n10667), .RESET_B(reset), .Q(n23800) );
  dfrtp_1 ___________________437785 ( .D(n10599), .CLK(n10666), .RESET_B(reset), .Q(n14) );
  dfrtp_1 ________________9_437610 ( .D(n10175), .CLK(n10658), .RESET_B(reset), 
        .Q(n23858) );
  dfrtp_1 ___________________437692 ( .D(n10182), .CLK(n10660), .RESET_B(reset), .Q(n23679) );
  dfrtp_1 ___________________437666 ( .D(n10181), .CLK(n10661), .RESET_B(reset), .Q(n23791) );
  dfrtp_1 ___________________437746 ( .D(n10180), .CLK(n10661), .RESET_B(reset), .Q(n13) );
  dfrtp_1 ___________________437688 ( .D(n10179), .CLK(n10661), .RESET_B(reset), .Q(n23790) );
  dfrtp_1 ___________________437400 ( .D(n10168), .CLK(n10664), .RESET_B(reset), .Q(n12) );
  dfrtp_1 ___________________437491 ( .D(n10169), .CLK(n10664), .RESET_B(reset), .Q(n23811) );
  dfrbp_1 ___________________437529 ( .D(n10548), .CLK(n10647), .RESET_B(reset), .Q_N(n755) );
  dfrtp_1 ___________________437552 ( .D(n10547), .CLK(n10664), .RESET_B(reset), .Q(n12478) );
  dfrtp_1 ___________________437417 ( .D(n10546), .CLK(n10664), .RESET_B(reset), .Q(n12442) );
  dfrtp_1 ___________________436916 ( .D(n10557), .CLK(n10666), .RESET_B(reset), .Q(n23909) );
  dfrtp_1 ___________________437347 ( .D(n10167), .CLK(n10664), .RESET_B(reset), .Q(n12581) );
  dfrtp_1 ___________________437381 ( .D(n10166), .CLK(n10656), .RESET_B(reset), .Q(n23826) );
  dfrtp_1 ___________________437430 ( .D(n10165), .CLK(n10664), .RESET_B(reset), .Q(n12582) );
  dfrtp_1 _________________9_437585 ( .D(n10183), .CLK(n10665), .RESET_B(reset), .Q(n23794) );
  dfrtp_1 ___________________437626 ( .D(n10214), .CLK(n10665), .RESET_B(reset), .Q(n23697) );
  dfrtp_1 ___________________437634 ( .D(n10215), .CLK(n10665), .RESET_B(reset), .Q(n23793) );
  dfrtp_1 ___________________437670 ( .D(n10184), .CLK(n10665), .RESET_B(reset), .Q(n12544) );
  dfrtp_1 _________________0_437231 ( .D(n10213), .CLK(n10666), .RESET_B(reset), .Q(n11) );
  dfrtp_1 ___________________437072 ( .D(n10436), .CLK(n10666), .RESET_B(reset), .Q(n12546) );
  dfrtp_1 ___________________437195 ( .D(n10174), .CLK(n10666), .RESET_B(reset), .Q(n10) );
  dfrtp_1 _________________9_437156 ( .D(n10437), .CLK(n10661), .RESET_B(reset), .Q(n9) );
  dfrtp_1 ___________________436979 ( .D(n10434), .CLK(n10661), .RESET_B(reset), .Q(n12515) );
  dfrtp_1 _________________0_437006 ( .D(n10433), .CLK(n10661), .RESET_B(reset), .Q(n8) );
  dfrbp_1 ___________________436915 ( .D(n10435), .CLK(n10648), .RESET_B(reset), .Q_N(n1519) );
  dfrbp_1 _________________9_437076 ( .D(n10432), .CLK(n10646), .RESET_B(reset), .Q(n10623), .Q_N(n1520) );
  dfrtp_1 ___________________436891 ( .D(n10569), .CLK(n10655), .RESET_B(reset), .Q(n7) );
  dfrtp_1 _____________9_____436735 ( .D(n10567), .CLK(n10655), .RESET_B(reset), .Q(n12511) );
  dfrtp_1 _________________0_436813 ( .D(n10530), .CLK(n10667), .RESET_B(reset), .Q(n23801) );
  dfrtp_1 ___________________437179 ( .D(n10171), .CLK(n10660), .RESET_B(reset), .Q(n23808) );
  dfrtp_1 ___________________437358 ( .D(n10170), .CLK(n10660), .RESET_B(reset), .Q(n23809) );
  dfrtp_1 ___________________437287 ( .D(n10173), .CLK(n10664), .RESET_B(reset), .Q(n12482) );
  dfrtp_1 ___________________437242 ( .D(n10172), .CLK(n10660), .RESET_B(reset), .Q(n6) );
  dfrbp_1 ___________________437057 ( .D(n10163), .CLK(n10646), .RESET_B(reset), .Q(n10644), .Q_N(n2113) );
  dfrtp_1 ___________________437180 ( .D(n10162), .CLK(n10664), .RESET_B(reset), .Q(n23702) );
  dfrbp_1 ___________________437129 ( .D(n10161), .CLK(n10649), .RESET_B(reset), .Q_N(n2116) );
  dfrtp_1 ___________________437050 ( .D(n10164), .CLK(n10664), .RESET_B(reset), .Q(n23676) );
  dfrtp_1 ___________________436653 ( .D(n10563), .CLK(n10652), .RESET_B(reset), .Q(n23941) );
  dfrtp_1 ___________________436770 ( .D(n10562), .CLK(n10661), .RESET_B(reset), .Q(n23942) );
  dfrtp_1 ___________________436876 ( .D(n10564), .CLK(n10655), .RESET_B(reset), .Q(n5) );
  dfrtp_1 _____________9___9_436427 ( .D(n10218), .CLK(n10660), .RESET_B(reset), .Q(n4) );
  dfrtp_1 ______________0_____436069 ( .D(n10429), .CLK(n10659), .RESET_B(
        reset), .Q(__________0_______18819) );
  dfrtp_1 ___________________436369 ( .D(n10431), .CLK(n10661), .RESET_B(reset), .Q(n23921) );
  dfrtp_1 _________________9_436553 ( .D(n10151), .CLK(n10658), .RESET_B(reset), .Q(n3) );
  dfrtp_1 _________________0_436533 ( .D(n10306), .CLK(n10668), .RESET_B(reset), .Q(n23705) );
  dfrtp_1 _________________0_ ( .D(n10590), .CLK(n10654), .RESET_B(reset), .Q(
        n2) );
  dfrtp_1 ___________________436493 ( .D(n10595), .CLK(n10668), .RESET_B(reset), .Q(_________________18785) );
  dfrtp_1 ___________________ ( .D(n10594), .CLK(n10668), .RESET_B(reset), .Q(
        n1) );
  dfrtp_1 _____________9_____ ( .D(n10593), .CLK(n10649), .RESET_B(reset), .Q(
        _________9_______18814) );
  inv_2 U10745 ( .A(n10677), .Y(n10648) );
  inv_2 U10746 ( .A(n10678), .Y(n10647) );
  inv_2 U10747 ( .A(n10675), .Y(n10649) );
  inv_2 U10748 ( .A(n10681), .Y(n10674) );
  inv_2 U10749 ( .A(n10680), .Y(n10670) );
  inv_2 U10750 ( .A(n10681), .Y(n10672) );
  inv_2 U10751 ( .A(n10680), .Y(n10671) );
  inv_2 U10752 ( .A(n10681), .Y(n10673) );
  inv_2 U10753 ( .A(n10675), .Y(n10653) );
  inv_2 U10754 ( .A(n10680), .Y(n10662) );
  inv_2 U10755 ( .A(n10679), .Y(n10666) );
  inv_2 U10756 ( .A(n10676), .Y(n10657) );
  inv_2 U10757 ( .A(n10676), .Y(n10656) );
  inv_2 U10758 ( .A(n10677), .Y(n10660) );
  inv_2 U10759 ( .A(n10675), .Y(n10652) );
  inv_2 U10760 ( .A(n10678), .Y(n10663) );
  inv_2 U10761 ( .A(n10679), .Y(n10667) );
  inv_2 U10762 ( .A(n10676), .Y(n10661) );
  inv_2 U10763 ( .A(n10681), .Y(n10651) );
  inv_2 U10764 ( .A(n10680), .Y(n10650) );
  inv_2 U10765 ( .A(n10678), .Y(n10665) );
  inv_2 U10766 ( .A(n10678), .Y(n10664) );
  inv_2 U10767 ( .A(n10679), .Y(n10668) );
  inv_2 U10768 ( .A(n10680), .Y(n10669) );
  inv_2 U10769 ( .A(n10676), .Y(n10655) );
  inv_2 U10770 ( .A(n10677), .Y(n10659) );
  inv_2 U10771 ( .A(n10675), .Y(n10654) );
  inv_2 U10772 ( .A(n10677), .Y(n10658) );
  inv_2 U10773 ( .A(n10679), .Y(n10646) );
  inv_2 U10774 ( .A(clk), .Y(n10681) );
  inv_2 U10775 ( .A(clk), .Y(n10678) );
  inv_2 U10776 ( .A(clk), .Y(n10679) );
  inv_2 U10777 ( .A(clk), .Y(n10680) );
  inv_2 U10778 ( .A(clk), .Y(n10676) );
  inv_2 U10779 ( .A(clk), .Y(n10675) );
  inv_2 U10780 ( .A(clk), .Y(n10677) );
  o21ai_0 U10781 ( .A1(n10682), .A2(n10683), .B1(n10684), .Y(n215) );
  mux2i_1 U10782 ( .A0(n10685), .A1(n10686), .S(n10687), .Y(n10684) );
  nor4_1 U10783 ( .A(n10688), .B(n10689), .C(n10690), .D(n10691), .Y(n10687)
         );
  nand3_1 U10784 ( .A(n10692), .B(n10693), .C(n10694), .Y(n10689) );
  nand4_1 U10785 ( .A(n10695), .B(n10696), .C(n10697), .D(n10698), .Y(n10688)
         );
  and3_1 U10786 ( .A(n10699), .B(n10700), .C(n10701), .X(n10698) );
  nor4_1 U10787 ( .A(n10702), .B(n10703), .C(n10704), .D(n10705), .Y(n10686)
         );
  nand2_1 U10788 ( .A(n10682), .B(n10706), .Y(n10703) );
  nand4_1 U10789 ( .A(n10707), .B(n10708), .C(n10709), .D(n10710), .Y(n10702)
         );
  and2_0 U10790 ( .A(n10711), .B(n10712), .X(n10682) );
  nor4_1 U10791 ( .A(n10713), .B(n10714), .C(n10715), .D(n10716), .Y(n10712)
         );
  inv_1 U10792 ( .A(n10717), .Y(n10714) );
  nand3_1 U10793 ( .A(n10718), .B(n10719), .C(n10720), .Y(n10713) );
  nor4_1 U10794 ( .A(n10721), .B(n10722), .C(n10723), .D(n10724), .Y(n10711)
         );
  nand3_1 U10795 ( .A(n10725), .B(n10726), .C(n10727), .Y(n10721) );
  o221ai_1 U10796 ( .A1(n10728), .A2(n10729), .B1(n10730), .B2(n10731), .C1(
        n10732), .Y(n209) );
  o21ai_0 U10797 ( .A1(n10733), .A2(n10734), .B1(n10735), .Y(n10732) );
  o21ai_0 U10798 ( .A1(n10736), .A2(n10737), .B1(n10738), .Y(n10734) );
  nor4_1 U10799 ( .A(n10739), .B(n10740), .C(n10741), .D(n10742), .Y(n10728)
         );
  nand3_1 U10800 ( .A(n10743), .B(n10744), .C(n10745), .Y(n10739) );
  o21ai_0 U10801 ( .A1(n10746), .A2(n10747), .B1(n10748), .Y(n198) );
  mux2i_1 U10802 ( .A0(n10749), .A1(n10750), .S(n10751), .Y(n10748) );
  nor4_1 U10803 ( .A(n10752), .B(n10753), .C(n10754), .D(n10755), .Y(n10751)
         );
  o21ai_0 U10804 ( .A1(n10756), .A2(n10757), .B1(n10758), .Y(n10753) );
  nand3_1 U10805 ( .A(n10759), .B(n10760), .C(n10761), .Y(n10752) );
  nor3_1 U10806 ( .A(n10762), .B(n10763), .C(n10764), .Y(n10750) );
  inv_1 U10807 ( .A(n10746), .Y(n10763) );
  nand3_1 U10808 ( .A(n10765), .B(n10697), .C(n10766), .Y(n10762) );
  nor4_1 U10809 ( .A(n10767), .B(n10768), .C(n10769), .D(n10770), .Y(n10746)
         );
  nand3_1 U10810 ( .A(n10771), .B(n10772), .C(n10773), .Y(n10770) );
  nor2_1 U10811 ( .A(n10774), .B(n10775), .Y(n10603) );
  nor2_1 U10812 ( .A(n10776), .B(n10774), .Y(n10602) );
  xor2_1 U10813 ( .A(n10777), .B(n10778), .X(n10776) );
  xnor2_1 U10814 ( .A(n23829), .B(n10779), .Y(n10778) );
  nand2_1 U10815 ( .A(n10780), .B(n10781), .Y(n10601) );
  mux2i_1 U10816 ( .A0(n10782), .A1(n10783), .S(n10784), .Y(n10780) );
  xnor2_1 U10817 ( .A(n10785), .B(n10786), .Y(n10783) );
  nand2_1 U10818 ( .A(n10787), .B(n10788), .Y(n10785) );
  inv_1 U10819 ( .A(n10789), .Y(n10787) );
  xor2_1 U10820 ( .A(n10635), .B(n10790), .X(n10782) );
  nand2_1 U10821 ( .A(n10791), .B(n10781), .Y(n10600) );
  mux2i_1 U10822 ( .A0(n10792), .A1(n10793), .S(n10784), .Y(n10791) );
  mux2i_1 U10823 ( .A0(n10794), .A1(n10795), .S(n10796), .Y(n10793) );
  nand2_1 U10824 ( .A(n10797), .B(n10798), .Y(n10795) );
  xnor2_1 U10825 ( .A(n10797), .B(n10798), .Y(n10794) );
  nand2_1 U10826 ( .A(inData[20]), .B(n10799), .Y(n10792) );
  xor2_1 U10827 ( .A(n10800), .B(n10790), .X(n10799) );
  nand2_1 U10828 ( .A(n31), .B(n10801), .Y(n10790) );
  inv_1 U10829 ( .A(n23840), .Y(n10801) );
  nor2_1 U10830 ( .A(n10802), .B(n10803), .Y(n10599) );
  xor2_1 U10831 ( .A(n10804), .B(n10805), .X(n10803) );
  xor2_1 U10832 ( .A(n10806), .B(n10807), .X(n10805) );
  xor2_1 U10833 ( .A(n10808), .B(n10809), .X(n10807) );
  o22ai_1 U10834 ( .A1(n10810), .A2(n10811), .B1(n10812), .B2(n10635), .Y(
        n10809) );
  nor2_1 U10835 ( .A(n23765), .B(n10813), .Y(n10812) );
  a21oi_1 U10836 ( .A1(n10814), .A2(n10815), .B1(n10816), .Y(n10806) );
  xor2_1 U10837 ( .A(n10817), .B(n10818), .X(n10804) );
  xor2_1 U10838 ( .A(n24045), .B(n12380), .X(n10818) );
  xor2_1 U10839 ( .A(n20745), .B(n31), .X(n10817) );
  o22ai_1 U10840 ( .A1(n10819), .A2(n10820), .B1(n10821), .B2(n10822), .Y(
        n10598) );
  xor2_1 U10841 ( .A(n23800), .B(n10823), .X(n10822) );
  xor2_1 U10842 ( .A(n10824), .B(n10825), .X(n10820) );
  xor2_1 U10843 ( .A(n10826), .B(n14), .X(n10825) );
  o22ai_1 U10844 ( .A1(n10827), .A2(n10828), .B1(n23680), .B2(n10829), .Y(
        n10824) );
  and2_0 U10845 ( .A(n10828), .B(n10827), .X(n10829) );
  o32ai_1 U10846 ( .A1(n10830), .A2(n10831), .A3(n10832), .B1(n10833), .B2(
        n10834), .Y(n10597) );
  xor2_1 U10847 ( .A(n10835), .B(n10836), .X(n10834) );
  xor2_1 U10848 ( .A(n10837), .B(n10838), .X(n10836) );
  xor2_1 U10849 ( .A(n10839), .B(n10840), .X(n10838) );
  o22ai_1 U10850 ( .A1(n10841), .A2(n10842), .B1(n10843), .B2(n10844), .Y(
        n10839) );
  and2_0 U10851 ( .A(n10842), .B(n10841), .X(n10843) );
  o22ai_1 U10852 ( .A1(n10827), .A2(n10845), .B1(n23721), .B2(n10846), .Y(
        n10837) );
  nor2_1 U10853 ( .A(n10847), .B(n10848), .Y(n10846) );
  xor2_1 U10854 ( .A(n12380), .B(n10849), .X(n10835) );
  xor2_1 U10855 ( .A(n66), .B(n23721), .X(n10849) );
  xor2_1 U10856 ( .A(n23882), .B(n23801), .X(n10830) );
  o22ai_1 U10857 ( .A1(n10832), .A2(n10850), .B1(n10851), .B2(n10833), .Y(
        n10596) );
  xor2_1 U10858 ( .A(n10852), .B(n10853), .X(n10851) );
  a21oi_1 U10859 ( .A1(n10854), .A2(n10855), .B1(n10856), .Y(n10853) );
  xor2_1 U10860 ( .A(n23885), .B(n23801), .X(n10850) );
  mux2i_1 U10861 ( .A0(n10857), .A1(n10858), .S(n10859), .Y(n10595) );
  xor2_1 U10862 ( .A(n10860), .B(n10861), .X(n10859) );
  o22ai_1 U10863 ( .A1(n10862), .A2(n10813), .B1(n23801), .B2(n10863), .Y(
        n10861) );
  and2_0 U10864 ( .A(n10813), .B(n10862), .X(n10863) );
  nand2_1 U10865 ( .A(n23922), .B(n10826), .Y(n10857) );
  nand2_1 U10866 ( .A(n23922), .B(n10864), .Y(n10594) );
  xor2_1 U10867 ( .A(n10865), .B(n10866), .X(n10864) );
  xor2_1 U10868 ( .A(n10867), .B(n10868), .X(n10866) );
  a21oi_1 U10869 ( .A1(n10869), .A2(n10870), .B1(n10871), .Y(n10867) );
  inv_1 U10870 ( .A(n10872), .Y(n10871) );
  or2_0 U10871 ( .A(n10873), .B(n10874), .X(n10870) );
  xor2_1 U10872 ( .A(n10875), .B(n10876), .X(n10865) );
  xor2_1 U10873 ( .A(n10877), .B(n10878), .X(n10876) );
  xor2_1 U10874 ( .A(n10879), .B(n10880), .X(n10878) );
  o22ai_1 U10875 ( .A1(n10881), .A2(n10882), .B1(n10883), .B2(n10884), .Y(
        n10880) );
  nor2_1 U10876 ( .A(n10885), .B(n10886), .Y(n10883) );
  inv_1 U10877 ( .A(n10882), .Y(n10885) );
  inv_1 U10878 ( .A(n10886), .Y(n10881) );
  xor2_1 U10879 ( .A(n10882), .B(n10887), .X(n10877) );
  a21oi_1 U10880 ( .A1(n10888), .A2(n12380), .B1(n10889), .Y(n10887) );
  a21oi_1 U10881 ( .A1(n10826), .A2(n10890), .B1(n23705), .Y(n10889) );
  inv_1 U10882 ( .A(n10888), .Y(n10890) );
  xor2_1 U10883 ( .A(n10891), .B(n10892), .X(n10875) );
  xor2_1 U10884 ( .A(outData[31]), .B(n23705), .X(n10892) );
  xor2_1 U10885 ( .A(n10893), .B(_________________18785), .X(n10891) );
  o32ai_1 U10886 ( .A1(n10894), .A2(n1), .A3(n10858), .B1(n10774), .B2(n10895), 
        .Y(n10593) );
  mux2i_1 U10887 ( .A0(n10896), .A1(n10897), .S(n1), .Y(n10895) );
  nand2_1 U10888 ( .A(n10898), .B(n10899), .Y(n10897) );
  inv_1 U10889 ( .A(n10900), .Y(n10899) );
  nand3_1 U10890 ( .A(n2), .B(n10826), .C(n10901), .Y(n10898) );
  inv_1 U10891 ( .A(n10902), .Y(n10896) );
  a21oi_1 U10892 ( .A1(n10894), .A2(n10901), .B1(n10903), .Y(n10902) );
  nand2_1 U10893 ( .A(n12380), .B(n23922), .Y(n10858) );
  inv_1 U10894 ( .A(n2), .Y(n10894) );
  nand2_1 U10895 ( .A(n23922), .B(n10904), .Y(n10592) );
  xor2_1 U10896 ( .A(n10905), .B(n10906), .X(n10904) );
  xor2_1 U10897 ( .A(n10882), .B(n10907), .X(n10906) );
  xor2_1 U10898 ( .A(n10908), .B(n10909), .X(n10907) );
  a21oi_1 U10899 ( .A1(n10910), .A2(n12318), .B1(n10911), .Y(n10909) );
  a21oi_1 U10900 ( .A1(n10912), .A2(n10913), .B1(n23898), .Y(n10911) );
  o22ai_1 U10901 ( .A1(n10914), .A2(n10915), .B1(n10916), .B2(n10884), .Y(
        n10908) );
  and2_0 U10902 ( .A(n10915), .B(n10914), .X(n10916) );
  xor2_1 U10903 ( .A(n10917), .B(n10918), .X(n10905) );
  xor2_1 U10904 ( .A(n10919), .B(n10920), .X(n10918) );
  xnor2_1 U10905 ( .A(n23898), .B(_________9_______18814), .Y(n10917) );
  o32ai_1 U10906 ( .A1(n10921), .A2(n10922), .A3(n10923), .B1(n23668), .B2(
        n10924), .Y(n10591) );
  xor2_1 U10907 ( .A(n23850), .B(n2046), .X(n10921) );
  nor2_1 U10908 ( .A(n10774), .B(n10925), .Y(n10590) );
  xor2_1 U10909 ( .A(n10869), .B(n10926), .X(n10925) );
  o21ai_0 U10910 ( .A1(n10874), .A2(n10873), .B1(n10872), .Y(n10926) );
  xor2_1 U10911 ( .A(n10927), .B(n10928), .X(n10872) );
  nand2_1 U10912 ( .A(n10874), .B(n10873), .Y(n10927) );
  xnor2_1 U10913 ( .A(n10884), .B(n10929), .Y(n10873) );
  xor2_1 U10914 ( .A(n10886), .B(n10882), .X(n10929) );
  xor2_1 U10915 ( .A(n10930), .B(n10931), .X(n10882) );
  xor2_1 U10916 ( .A(outData[31]), .B(n10932), .X(n10931) );
  nor2_1 U10917 ( .A(n10933), .B(n10934), .Y(n10932) );
  xor2_1 U10918 ( .A(n10935), .B(n10936), .X(n10934) );
  nand2_1 U10919 ( .A(n10937), .B(n10938), .Y(n10935) );
  inv_1 U10920 ( .A(n10939), .Y(n10933) );
  nand2_1 U10921 ( .A(n10940), .B(n10941), .Y(n10886) );
  xor2_1 U10922 ( .A(n10942), .B(n10943), .X(n10941) );
  nor2_1 U10923 ( .A(n10944), .B(n10945), .Y(n10943) );
  xor2_1 U10924 ( .A(n10946), .B(n10947), .X(n10940) );
  nor2_1 U10925 ( .A(n10948), .B(n10949), .Y(n10947) );
  xnor2_1 U10926 ( .A(n10888), .B(n10950), .Y(n10874) );
  xor2_1 U10927 ( .A(n23705), .B(n12380), .X(n10950) );
  a22oi_1 U10928 ( .A1(n10810), .A2(n10951), .B1(n10952), .B2(n3), .Y(n10888)
         );
  or2_0 U10929 ( .A(n10951), .B(n10810), .X(n10952) );
  o21ai_0 U10930 ( .A1(n10953), .A2(n10954), .B1(n10955), .Y(n10869) );
  xor2_1 U10931 ( .A(n10808), .B(n10956), .X(n10955) );
  nand2_1 U10932 ( .A(n23922), .B(n10957), .Y(n10589) );
  xor2_1 U10933 ( .A(n10958), .B(n10959), .X(n10957) );
  nor2_1 U10934 ( .A(n10900), .B(n10960), .Y(n10959) );
  mux2i_1 U10935 ( .A0(n10961), .A1(n10962), .S(n2), .Y(n10960) );
  a21oi_1 U10936 ( .A1(n10901), .A2(n12380), .B1(n10903), .Y(n10962) );
  nor3_1 U10937 ( .A(n10901), .B(n2), .C(n10826), .Y(n10900) );
  a21oi_1 U10938 ( .A1(n10963), .A2(n23934), .B1(n10903), .Y(n10901) );
  a21oi_1 U10939 ( .A1(n10964), .A2(n10965), .B1(n12380), .Y(n10903) );
  nor2_1 U10940 ( .A(n10774), .B(n10966), .Y(n10588) );
  xnor2_1 U10941 ( .A(n10914), .B(n10967), .Y(n10966) );
  xor2_1 U10942 ( .A(n10915), .B(n10884), .X(n10967) );
  o22ai_1 U10943 ( .A1(n10968), .A2(n10969), .B1(n10970), .B2(n10971), .Y(
        n10915) );
  and2_0 U10944 ( .A(n10969), .B(n10968), .X(n10971) );
  xor2_1 U10945 ( .A(n10972), .B(n10973), .X(n10914) );
  xor2_1 U10946 ( .A(n23903), .B(n23898), .X(n10973) );
  xor2_1 U10947 ( .A(n10912), .B(n10910), .X(n10972) );
  inv_1 U10948 ( .A(n10913), .Y(n10910) );
  o22ai_1 U10949 ( .A1(n10974), .A2(n10912), .B1(n10975), .B2(n10629), .Y(
        n10913) );
  and2_0 U10950 ( .A(n10974), .B(n10912), .X(n10975) );
  inv_1 U10951 ( .A(n12318), .Y(n10912) );
  o211ai_1 U10952 ( .A1(n10976), .A2(n10977), .B1(n10978), .C1(n10979), .Y(
        n10587) );
  mux2i_1 U10953 ( .A0(n10980), .A1(n10981), .S(n10982), .Y(n10979) );
  nor4_1 U10954 ( .A(n10983), .B(n10984), .C(n10985), .D(n10986), .Y(n10982)
         );
  o21ai_0 U10955 ( .A1(n10987), .A2(n10988), .B1(n10989), .Y(n10984) );
  nand4_1 U10956 ( .A(n10990), .B(n10991), .C(n10992), .D(n10993), .Y(n10983)
         );
  and2_0 U10957 ( .A(n10994), .B(n10995), .X(n10993) );
  nor4_1 U10958 ( .A(n10996), .B(n10997), .C(n10998), .D(n10999), .Y(n10981)
         );
  nand2_1 U10959 ( .A(n11000), .B(n11001), .Y(n10999) );
  nand3_1 U10960 ( .A(n11002), .B(n11003), .C(n11004), .Y(n10997) );
  nand4_1 U10961 ( .A(n11005), .B(n11006), .C(n11007), .D(n11008), .Y(n10996)
         );
  nor4_1 U10962 ( .A(n11009), .B(n11010), .C(n11011), .D(n11012), .Y(n11008)
         );
  inv_1 U10963 ( .A(n11013), .Y(n10976) );
  o21ai_0 U10964 ( .A1(n11014), .A2(n11005), .B1(n11002), .Y(n11013) );
  and4_1 U10965 ( .A(n11015), .B(n11016), .C(n11017), .D(n11018), .X(n11002)
         );
  nor4_1 U10966 ( .A(n11019), .B(n11020), .C(n11021), .D(n11022), .Y(n11018)
         );
  inv_1 U10967 ( .A(n11023), .Y(n11022) );
  nand3_1 U10968 ( .A(n11024), .B(n11025), .C(n11026), .Y(n11019) );
  nor3_1 U10969 ( .A(n11027), .B(n11028), .C(n11029), .Y(n11017) );
  inv_1 U10970 ( .A(n11030), .Y(n11028) );
  nand2_1 U10971 ( .A(n11031), .B(n11032), .Y(n10586) );
  mux2i_1 U10972 ( .A0(n11033), .A1(n11034), .S(n11035), .Y(n11031) );
  nand2_1 U10973 ( .A(n11036), .B(inData[14]), .Y(n11034) );
  xor2_1 U10974 ( .A(n11037), .B(n20), .X(n11036) );
  nand2_1 U10975 ( .A(n23878), .B(n23877), .Y(n11037) );
  xor2_1 U10976 ( .A(n11038), .B(n11039), .X(n11033) );
  a21oi_1 U10977 ( .A1(n11040), .A2(n11041), .B1(n11042), .Y(n11038) );
  mux2i_1 U10978 ( .A0(n11043), .A1(n11044), .S(n11035), .Y(n10585) );
  nand2_1 U10979 ( .A(n11045), .B(n11046), .Y(n11044) );
  xor2_1 U10980 ( .A(n11047), .B(n11048), .X(n11043) );
  xnor2_1 U10981 ( .A(n11049), .B(n11050), .Y(n11047) );
  nor2_1 U10982 ( .A(n11051), .B(n11052), .Y(n11050) );
  nand2_1 U10983 ( .A(n11053), .B(n11032), .Y(n10584) );
  mux2i_1 U10984 ( .A0(n11054), .A1(n11055), .S(n11035), .Y(n11053) );
  nand2_1 U10985 ( .A(inData[10]), .B(n23878), .Y(n11055) );
  xor2_1 U10986 ( .A(n11056), .B(n23979), .X(n11054) );
  o32ai_1 U10987 ( .A1(n11057), .A2(n11058), .A3(n11059), .B1(n11060), .B2(
        n11061), .Y(n11056) );
  nor2_1 U10988 ( .A(n11062), .B(n11063), .Y(n11060) );
  inv_1 U10989 ( .A(n11064), .Y(n11059) );
  o21ai_0 U10990 ( .A1(n11063), .A2(n11062), .B1(n11065), .Y(n11064) );
  o32ai_1 U10991 ( .A1(n11066), .A2(n10831), .A3(n10630), .B1(n11067), .B2(
        n11068), .Y(n10583) );
  xor2_1 U10992 ( .A(n11069), .B(n11070), .X(n11067) );
  xor2_1 U10993 ( .A(n23877), .B(n11071), .X(n11069) );
  mux2i_1 U10994 ( .A0(n11072), .A1(n11073), .S(n11068), .Y(n10582) );
  a211oi_1 U10995 ( .A1(n11074), .A2(n11075), .B1(n11076), .C1(n11077), .Y(
        n11073) );
  inv_1 U10996 ( .A(n11078), .Y(n11077) );
  o21ai_0 U10997 ( .A1(n20747), .A2(n41), .B1(inData[8]), .Y(n11076) );
  a21oi_1 U10998 ( .A1(n11079), .A2(n11080), .B1(n11081), .Y(n11072) );
  a21oi_1 U10999 ( .A1(n11082), .A2(n11080), .B1(n11083), .Y(n11081) );
  o32ai_1 U11000 ( .A1(n11084), .A2(n11085), .A3(n11086), .B1(n11087), .B2(
        n11088), .Y(n10581) );
  xnor2_1 U11001 ( .A(n11089), .B(n11090), .Y(n11088) );
  xor2_1 U11002 ( .A(n11091), .B(n11092), .X(n11090) );
  xor2_1 U11003 ( .A(n11093), .B(n23687), .X(n11085) );
  nand2_1 U11004 ( .A(n23861), .B(n23786), .Y(n11093) );
  o32ai_1 U11005 ( .A1(n11094), .A2(n11095), .A3(n10923), .B1(n11096), .B2(
        n11097), .Y(n10580) );
  xor2_1 U11006 ( .A(n11098), .B(n11099), .X(n11096) );
  xor2_1 U11007 ( .A(n11100), .B(n11101), .X(n11099) );
  xor2_1 U11008 ( .A(n11102), .B(n11103), .X(n11098) );
  xor2_1 U11009 ( .A(n11104), .B(n23786), .X(n11095) );
  nand2_1 U11010 ( .A(n23861), .B(n11105), .Y(n11104) );
  o32ai_1 U11011 ( .A1(n11094), .A2(n11106), .A3(n11107), .B1(n11097), .B2(
        n11108), .Y(n10579) );
  xor2_1 U11012 ( .A(n11109), .B(n11110), .X(n11108) );
  nand2_1 U11013 ( .A(n11111), .B(n11112), .Y(n11110) );
  nand2_1 U11014 ( .A(n11113), .B(n11114), .Y(n10578) );
  mux2i_1 U11015 ( .A0(n11115), .A1(n11116), .S(n11117), .Y(n11113) );
  o21ai_0 U11016 ( .A1(n20748), .A2(n11118), .B1(n11119), .Y(n11116) );
  xor2_1 U11017 ( .A(n11120), .B(n11121), .X(n11115) );
  xor2_1 U11018 ( .A(n23861), .B(n11122), .X(n11121) );
  nand2_1 U11019 ( .A(n11123), .B(n11114), .Y(n10577) );
  mux2i_1 U11020 ( .A0(n11124), .A1(n11125), .S(n11117), .Y(n11123) );
  nand2_1 U11021 ( .A(n11126), .B(n10646), .Y(n11125) );
  xor2_1 U11022 ( .A(n11119), .B(n23869), .X(n11126) );
  xor2_1 U11023 ( .A(n11127), .B(n11128), .X(n11124) );
  xor2_1 U11024 ( .A(n11129), .B(n11130), .X(n11128) );
  xor2_1 U11025 ( .A(n10628), .B(n11131), .X(n11127) );
  o32ai_1 U11026 ( .A1(n11132), .A2(n11133), .A3(n11134), .B1(n11117), .B2(
        n11135), .Y(n10576) );
  xor2_1 U11027 ( .A(n11136), .B(n11137), .X(n11135) );
  xor2_1 U11028 ( .A(n11138), .B(n23712), .X(n11137) );
  xnor2_1 U11029 ( .A(n23864), .B(n11119), .Y(n11132) );
  nand2_1 U11030 ( .A(n20748), .B(n11118), .Y(n11119) );
  mux2i_1 U11031 ( .A0(n11139), .A1(n11140), .S(n11141), .Y(n10575) );
  xor2_1 U11032 ( .A(n11142), .B(n11143), .X(n11140) );
  xor2_1 U11033 ( .A(n11144), .B(n11145), .X(n11143) );
  xor2_1 U11034 ( .A(n10936), .B(n11146), .X(n11142) );
  nand3_1 U11035 ( .A(n11147), .B(n11148), .C(inData[2]), .Y(n11139) );
  xor2_1 U11036 ( .A(n54), .B(n23969), .X(n11147) );
  o22ai_1 U11037 ( .A1(n11149), .A2(n11150), .B1(n11151), .B2(n11152), .Y(
        n10574) );
  xor2_1 U11038 ( .A(n11153), .B(n11154), .X(n11151) );
  a21oi_1 U11039 ( .A1(n12473), .A2(n11155), .B1(n11156), .Y(n11154) );
  nand2_1 U11040 ( .A(n23922), .B(n11157), .Y(n10573) );
  xor2_1 U11041 ( .A(n11158), .B(n11159), .X(n11157) );
  o22ai_1 U11042 ( .A1(n11160), .A2(n11161), .B1(n11162), .B2(n11163), .Y(
        n11158) );
  a21oi_1 U11043 ( .A1(n11164), .A2(n11165), .B1(n11160), .Y(n11162) );
  mux2_1 U11044 ( .A0(n11166), .A1(n11167), .S(n11165), .X(n11161) );
  nor3_1 U11045 ( .A(n11168), .B(n11164), .C(n11165), .Y(n11160) );
  mux2_1 U11046 ( .A0(______9__34498), .A1(n11169), .S(n11170), .X(n10572) );
  nand2_1 U11047 ( .A(n11171), .B(n11172), .Y(n11169) );
  xor2_1 U11048 ( .A(outData[14]), .B(n11173), .X(n11172) );
  inv_1 U11049 ( .A(n11174), .Y(n11171) );
  o32ai_1 U11050 ( .A1(n11175), .A2(n11176), .A3(n11177), .B1(n23666), .B2(
        n11170), .Y(n10571) );
  xor2_1 U11051 ( .A(n10611), .B(n11173), .X(n11176) );
  nand3_1 U11052 ( .A(n11178), .B(n11179), .C(n11180), .Y(n10570) );
  mux2i_1 U11053 ( .A0(n11181), .A1(n11182), .S(n11141), .Y(n11180) );
  xor2_1 U11054 ( .A(n11183), .B(n11184), .X(n11182) );
  xor2_1 U11055 ( .A(n11185), .B(n11186), .X(n11184) );
  xor2_1 U11056 ( .A(n11187), .B(n11188), .X(n11183) );
  and2_0 U11057 ( .A(n23909), .B(n23945), .X(n11181) );
  o211ai_1 U11058 ( .A1(n23946), .A2(n11179), .B1(n11178), .C1(n11189), .Y(
        n10569) );
  mux2i_1 U11059 ( .A0(n11190), .A1(n11191), .S(n11141), .Y(n11189) );
  xnor2_1 U11060 ( .A(n11192), .B(n11193), .Y(n11191) );
  xor2_1 U11061 ( .A(n11194), .B(n11195), .X(n11192) );
  o21ai_0 U11062 ( .A1(n11196), .A2(n11197), .B1(inData[20]), .Y(n11190) );
  o211ai_1 U11063 ( .A1(n11198), .A2(n11199), .B1(n11178), .C1(n11200), .Y(
        n10568) );
  mux2i_1 U11064 ( .A0(n11201), .A1(n11202), .S(n7), .Y(n11200) );
  nor2_1 U11065 ( .A(n11141), .B(n11196), .Y(n11202) );
  inv_1 U11066 ( .A(n11179), .Y(n11201) );
  nand2_1 U11067 ( .A(n11196), .B(n11199), .Y(n11179) );
  nor2_1 U11068 ( .A(n23945), .B(n23909), .Y(n11196) );
  inv_1 U11069 ( .A(n11141), .Y(n11199) );
  xor2_1 U11070 ( .A(n11203), .B(n11204), .X(n11198) );
  xor2_1 U11071 ( .A(n11205), .B(n11206), .X(n11204) );
  nand2_1 U11072 ( .A(n11207), .B(n11208), .Y(n11203) );
  xor2_1 U11073 ( .A(n11209), .B(n11210), .X(n11207) );
  o32ai_1 U11074 ( .A1(n11211), .A2(n11212), .A3(n10923), .B1(n11213), .B2(
        n11214), .Y(n10567) );
  xnor2_1 U11075 ( .A(n7), .B(n11215), .Y(n11214) );
  nand2_1 U11076 ( .A(n11216), .B(n11217), .Y(n11215) );
  inv_1 U11077 ( .A(n11218), .Y(n11216) );
  nor2_1 U11078 ( .A(n11219), .B(n10774), .Y(n10566) );
  xnor2_1 U11079 ( .A(n11220), .B(n11221), .Y(n11219) );
  xor2_1 U11080 ( .A(n11222), .B(n11223), .X(n11221) );
  mux2i_1 U11081 ( .A0(n29), .A1(n11224), .S(n11170), .Y(n10565) );
  nor2_1 U11082 ( .A(n11225), .B(n11226), .Y(n11224) );
  nand2_1 U11083 ( .A(n11227), .B(n11228), .Y(n10564) );
  mux2i_1 U11084 ( .A0(n11229), .A1(n11230), .S(n11231), .Y(n11227) );
  xnor2_1 U11085 ( .A(n11232), .B(n11233), .Y(n11230) );
  xor2_1 U11086 ( .A(n11234), .B(n11235), .X(n11233) );
  nand2_1 U11087 ( .A(n11236), .B(inData[22]), .Y(n11229) );
  xor2_1 U11088 ( .A(n11237), .B(n23943), .X(n11236) );
  nand2_1 U11089 ( .A(n11238), .B(n11228), .Y(n10563) );
  mux2i_1 U11090 ( .A0(n11239), .A1(n11240), .S(n11231), .Y(n11238) );
  o22ai_1 U11091 ( .A1(n11241), .A2(n11242), .B1(n11243), .B2(n11244), .Y(
        n11240) );
  nor2_1 U11092 ( .A(n11241), .B(n11245), .Y(n11243) );
  inv_1 U11093 ( .A(n11246), .Y(n11242) );
  xor2_1 U11094 ( .A(n11247), .B(n11248), .X(n11239) );
  xor2_1 U11095 ( .A(n5), .B(n23942), .X(n11248) );
  nand2_1 U11096 ( .A(n23943), .B(n11249), .Y(n11247) );
  nand2_1 U11097 ( .A(n11250), .B(n11228), .Y(n10562) );
  mux2i_1 U11098 ( .A0(n23941), .A1(n11251), .S(n11231), .Y(n11250) );
  xor2_1 U11099 ( .A(n11252), .B(n11253), .X(n11251) );
  o21ai_0 U11100 ( .A1(n11254), .A2(n11255), .B1(n11256), .Y(n11253) );
  mux2i_1 U11101 ( .A0(n11257), .A1(n11258), .S(n11231), .Y(n10561) );
  xor2_1 U11102 ( .A(n11259), .B(n11260), .X(n11258) );
  nand2_1 U11103 ( .A(n11261), .B(n11262), .Y(n11259) );
  nand3_1 U11104 ( .A(n11263), .B(n11237), .C(inData[24]), .Y(n11257) );
  o21ai_0 U11105 ( .A1(n11213), .A2(n11264), .B1(n11265), .Y(n10560) );
  mux2i_1 U11106 ( .A0(n11266), .A1(n11267), .S(n62), .Y(n11265) );
  xor2_1 U11107 ( .A(n11268), .B(n11269), .X(n11264) );
  nand2_1 U11108 ( .A(n11270), .B(n11271), .Y(n11269) );
  nand2_1 U11109 ( .A(n23922), .B(n11272), .Y(n10559) );
  xnor2_1 U11110 ( .A(n11273), .B(n11274), .Y(n11272) );
  nand2_1 U11111 ( .A(n11275), .B(n11276), .Y(n11273) );
  o22ai_1 U11112 ( .A1(n57), .A2(n11170), .B1(n11277), .B2(n11177), .Y(n10558)
         );
  xor2_1 U11113 ( .A(outData[16]), .B(n12346), .X(n11277) );
  nand2_1 U11114 ( .A(n11278), .B(n11178), .Y(n10557) );
  mux2i_1 U11115 ( .A0(n23945), .A1(n11279), .S(n11141), .Y(n11278) );
  xor2_1 U11116 ( .A(n11280), .B(n11281), .X(n11279) );
  xor2_1 U11117 ( .A(n11282), .B(n11283), .X(n11281) );
  xor2_1 U11118 ( .A(n11284), .B(n11285), .X(n11280) );
  mux2i_1 U11119 ( .A0(n11286), .A1(n11287), .S(n11213), .Y(n10556) );
  a211oi_1 U11120 ( .A1(n11212), .A2(n11288), .B1(n11289), .C1(n11134), .Y(
        n11287) );
  xor2_1 U11121 ( .A(n11290), .B(n11291), .X(n11286) );
  xnor2_1 U11122 ( .A(n11292), .B(n11293), .Y(n11291) );
  xor2_1 U11123 ( .A(n23945), .B(n11294), .X(n11293) );
  xor2_1 U11124 ( .A(n11295), .B(n11296), .X(n11290) );
  nor2_1 U11125 ( .A(n10774), .B(n11297), .Y(n10555) );
  xor2_1 U11126 ( .A(n11298), .B(n11299), .X(n11297) );
  xor2_1 U11127 ( .A(n11300), .B(n11301), .X(n11299) );
  nand2_1 U11128 ( .A(n11302), .B(n11303), .Y(n11298) );
  o21ai_0 U11129 ( .A1(n12413), .A2(n11304), .B1(n11305), .Y(n10554) );
  nand2_1 U11130 ( .A(__________0_____), .B(n11306), .Y(n11305) );
  nand2_1 U11131 ( .A(n11307), .B(n11178), .Y(n10553) );
  or2_0 U11132 ( .A(n11148), .B(n11141), .X(n11178) );
  nand4_1 U11133 ( .A(n11308), .B(n11309), .C(n11310), .D(n11311), .Y(n11148)
         );
  mux2i_1 U11134 ( .A0(n11312), .A1(n11313), .S(n11141), .Y(n11307) );
  a211oi_1 U11135 ( .A1(n11314), .A2(n11315), .B1(n11316), .C1(n11317), .Y(
        n11141) );
  o221ai_1 U11136 ( .A1(n11318), .A2(n11319), .B1(n11311), .B2(n11320), .C1(
        n11321), .Y(n11317) );
  o22ai_1 U11137 ( .A1(n11322), .A2(n11323), .B1(n11324), .B2(n11325), .Y(
        n11313) );
  a21oi_1 U11138 ( .A1(n11326), .A2(n11327), .B1(n11322), .Y(n11324) );
  inv_1 U11139 ( .A(n11328), .Y(n11323) );
  xor2_1 U11140 ( .A(n11329), .B(n12473), .X(n11312) );
  nand2_1 U11141 ( .A(n54), .B(n698), .Y(n11329) );
  o32ai_1 U11142 ( .A1(n11330), .A2(n10638), .A3(n11331), .B1(n11332), .B2(
        n11333), .Y(n10552) );
  xor2_1 U11143 ( .A(n11334), .B(n11335), .X(n11332) );
  xor2_1 U11144 ( .A(n11336), .B(n11337), .X(n11335) );
  o21ai_0 U11145 ( .A1(n11338), .A2(n11339), .B1(n11340), .Y(n11334) );
  o22ai_1 U11146 ( .A1(n11341), .A2(n11152), .B1(n11342), .B2(n11150), .Y(
        n10551) );
  xor2_1 U11147 ( .A(n11343), .B(n49), .X(n11342) );
  xor2_1 U11148 ( .A(n11344), .B(n11345), .X(n11341) );
  xor2_1 U11149 ( .A(n54), .B(n11346), .X(n11345) );
  xor2_1 U11150 ( .A(n11347), .B(n11348), .X(n11344) );
  nand2_1 U11151 ( .A(n11349), .B(n23922), .Y(n10550) );
  xor2_1 U11152 ( .A(n11350), .B(n11351), .X(n11349) );
  nor2_1 U11153 ( .A(n11352), .B(n11353), .Y(n11351) );
  inv_1 U11154 ( .A(n11354), .Y(n11352) );
  o32ai_1 U11155 ( .A1(n11355), .A2(n11304), .A3(n11356), .B1(n23669), .B2(
        n11357), .Y(n10549) );
  xor2_1 U11156 ( .A(outData[9]), .B(n12330), .X(n11356) );
  mux2i_1 U11157 ( .A0(n11358), .A1(n11359), .S(n11360), .Y(n10548) );
  xnor2_1 U11158 ( .A(n11361), .B(n11362), .Y(n11359) );
  nand2_1 U11159 ( .A(n11363), .B(n11364), .Y(n11361) );
  nor2_1 U11160 ( .A(n11365), .B(n11366), .Y(n11358) );
  o32ai_1 U11161 ( .A1(n11367), .A2(n11368), .A3(n11369), .B1(n11370), .B2(
        n11371), .Y(n10547) );
  xor2_1 U11162 ( .A(n11372), .B(n11373), .X(n11371) );
  xnor2_1 U11163 ( .A(n11374), .B(n11375), .Y(n11373) );
  xor2_1 U11164 ( .A(n11376), .B(n23995), .X(n11372) );
  xor2_1 U11165 ( .A(n11365), .B(n755), .X(n11369) );
  nand3_1 U11166 ( .A(n11377), .B(n11378), .C(n11379), .Y(n10546) );
  mux2i_1 U11167 ( .A0(n11380), .A1(n11381), .S(n11382), .Y(n11379) );
  xor2_1 U11168 ( .A(n11383), .B(n11384), .X(n11381) );
  xor2_1 U11169 ( .A(n24045), .B(n12478), .X(n11384) );
  xor2_1 U11170 ( .A(n11385), .B(n11386), .X(n11383) );
  o21ai_0 U11171 ( .A1(n11387), .A2(n11388), .B1(inData[10]), .Y(n11380) );
  inv_1 U11172 ( .A(n23826), .Y(n11387) );
  nand2_1 U11173 ( .A(n11389), .B(n11390), .Y(n10545) );
  mux2i_1 U11174 ( .A0(n11391), .A1(n11392), .S(n11393), .Y(n11389) );
  o21ai_0 U11175 ( .A1(n23704), .A2(n11394), .B1(n11395), .Y(n11392) );
  xor2_1 U11176 ( .A(n11396), .B(n11397), .X(n11391) );
  xor2_1 U11177 ( .A(n11398), .B(n11399), .X(n11396) );
  o32ai_1 U11178 ( .A1(n11107), .A2(n68), .A3(n11400), .B1(n11401), .B2(n11402), .Y(n10544) );
  xnor2_1 U11179 ( .A(n11403), .B(n11404), .Y(n11401) );
  xor2_1 U11180 ( .A(n756), .B(n11405), .X(n11403) );
  nor2_1 U11181 ( .A(n10774), .B(n11406), .Y(n10543) );
  xor2_1 U11182 ( .A(n11407), .B(n11408), .X(n11406) );
  xnor2_1 U11183 ( .A(n11409), .B(n11410), .Y(n11408) );
  xnor2_1 U11184 ( .A(n11411), .B(n11412), .Y(n11407) );
  xor2_1 U11185 ( .A(n11413), .B(n11414), .X(n11412) );
  o21ai_0 U11186 ( .A1(n11415), .A2(n11416), .B1(n11417), .Y(n10542) );
  nand2_1 U11187 ( .A(__________0_______18820), .B(n11418), .Y(n11417) );
  o21ai_0 U11188 ( .A1(n11419), .A2(n11420), .B1(n11421), .Y(n10541) );
  nand2_1 U11189 ( .A(n23870), .B(n11418), .Y(n11421) );
  xor2_1 U11190 ( .A(n11422), .B(outData[26]), .X(n11419) );
  nand2_1 U11191 ( .A(outData[24]), .B(outData[25]), .Y(n11422) );
  nand2_1 U11192 ( .A(n11423), .B(n11228), .Y(n10540) );
  or2_0 U11193 ( .A(n11263), .B(n11231), .X(n11228) );
  mux2i_1 U11194 ( .A0(n11424), .A1(n11425), .S(n11231), .Y(n11423) );
  xor2_1 U11195 ( .A(n11426), .B(n11427), .X(n11425) );
  xor2_1 U11196 ( .A(n11292), .B(n11428), .X(n11427) );
  o22ai_1 U11197 ( .A1(n11429), .A2(n11430), .B1(n11431), .B2(n11432), .Y(
        n11426) );
  nor2_1 U11198 ( .A(n11433), .B(n11429), .Y(n11431) );
  nand2_1 U11199 ( .A(inData[20]), .B(n11394), .Y(n11424) );
  mux2i_1 U11200 ( .A0(n11434), .A1(n11435), .S(n11231), .Y(n10539) );
  and4_1 U11201 ( .A(n11321), .B(n11309), .C(n11436), .D(n11437), .X(n11231)
         );
  a211oi_1 U11202 ( .A1(n11438), .A2(n24061), .B1(n11439), .C1(n11440), .Y(
        n11437) );
  a21oi_1 U11203 ( .A1(n11319), .A2(n11441), .B1(n11442), .Y(n11440) );
  nor3_1 U11204 ( .A(n11443), .B(n11444), .C(n11445), .Y(n11439) );
  xor2_1 U11205 ( .A(n11446), .B(n11447), .X(n11435) );
  xor2_1 U11206 ( .A(n11448), .B(n11449), .X(n11447) );
  nand2_1 U11207 ( .A(n11450), .B(n11263), .Y(n11434) );
  nand3_1 U11208 ( .A(n11318), .B(n11451), .C(n11452), .Y(n11263) );
  a22oi_1 U11209 ( .A1(n11453), .A2(n11315), .B1(n24061), .B2(n11454), .Y(
        n11452) );
  o21ai_0 U11210 ( .A1(n11394), .A2(n10633), .B1(n11395), .Y(n11450) );
  mux2_1 U11211 ( .A0(n10633), .A1(n11455), .S(n23704), .X(n11395) );
  nand2_1 U11212 ( .A(n10633), .B(n11394), .Y(n11455) );
  o22ai_1 U11213 ( .A1(n11400), .A2(n11456), .B1(n11457), .B2(n11402), .Y(
        n10538) );
  xor2_1 U11214 ( .A(n11458), .B(n11459), .X(n11457) );
  xnor2_1 U11215 ( .A(n23704), .B(n11460), .Y(n11459) );
  xor2_1 U11216 ( .A(n4), .B(n11461), .X(n11456) );
  nand2_1 U11217 ( .A(n11462), .B(n23922), .Y(n10537) );
  xor2_1 U11218 ( .A(n11463), .B(n11464), .X(n11462) );
  mux2i_1 U11219 ( .A0(n11465), .A1(n11466), .S(n11467), .Y(n11463) );
  o32ai_1 U11220 ( .A1(n11355), .A2(n12426), .A3(n11415), .B1(_____9___34413), 
        .B2(n10924), .Y(n10536) );
  o21ai_0 U11221 ( .A1(n11415), .A2(n11468), .B1(n11469), .Y(n10535) );
  nand2_1 U11222 ( .A(__________0___0___18817), .B(n11418), .Y(n11469) );
  o22ai_1 U11223 ( .A1(n11470), .A2(n11471), .B1(n11472), .B2(n11473), .Y(
        n10534) );
  o21ai_0 U11224 ( .A1(n23997), .A2(n821), .B1(n11474), .Y(n11473) );
  xnor2_1 U11225 ( .A(n11475), .B(n11476), .Y(n11471) );
  nor2_1 U11226 ( .A(n11477), .B(n11478), .Y(n11476) );
  inv_1 U11227 ( .A(n11479), .Y(n11477) );
  o32ai_1 U11228 ( .A1(n11480), .A2(n12467), .A3(n11134), .B1(n11481), .B2(
        n11482), .Y(n10533) );
  xor2_1 U11229 ( .A(n11483), .B(n11484), .X(n11481) );
  xor2_1 U11230 ( .A(n11485), .B(n23936), .X(n11483) );
  nand2_1 U11231 ( .A(n23922), .B(n11486), .Y(n10532) );
  xor2_1 U11232 ( .A(n11487), .B(n11488), .X(n11486) );
  xor2_1 U11233 ( .A(n11489), .B(n11490), .X(n11488) );
  nor2_1 U11234 ( .A(n11491), .B(n11492), .Y(n11487) );
  inv_1 U11235 ( .A(n11493), .Y(n11491) );
  mux2_1 U11236 ( .A0(n11494), .A1(______0__34499), .S(n11418), .X(n10531) );
  nand4_1 U11237 ( .A(inData[14]), .B(n11495), .C(n11496), .D(n11497), .Y(
        n11494) );
  nand2_1 U11238 ( .A(n10612), .B(n11498), .Y(n11496) );
  nand2_1 U11239 ( .A(n11499), .B(n11500), .Y(n10530) );
  mux2i_1 U11240 ( .A0(n11501), .A1(n11502), .S(n11503), .Y(n11499) );
  xor2_1 U11241 ( .A(n10844), .B(n11504), .X(n11502) );
  xor2_1 U11242 ( .A(n10841), .B(n10842), .X(n11504) );
  xnor2_1 U11243 ( .A(n10848), .B(n11505), .Y(n10842) );
  xor2_1 U11244 ( .A(n23721), .B(n10847), .X(n11505) );
  inv_1 U11245 ( .A(n11506), .Y(n10841) );
  o21ai_0 U11246 ( .A1(n11507), .A2(n11508), .B1(n11509), .Y(n11506) );
  xor2_1 U11247 ( .A(n11510), .B(n11511), .X(n11507) );
  xor2_1 U11248 ( .A(n11512), .B(n23903), .X(n10844) );
  o22ai_1 U11249 ( .A1(n11513), .A2(n11514), .B1(n10856), .B2(n10852), .Y(
        n11512) );
  o22ai_1 U11250 ( .A1(n11515), .A2(n11516), .B1(n11517), .B2(n11518), .Y(
        n10852) );
  inv_1 U11251 ( .A(n11519), .Y(n11518) );
  and2_0 U11252 ( .A(n11516), .B(n11515), .X(n11517) );
  xor2_1 U11253 ( .A(n11520), .B(n11521), .X(n10856) );
  nor2_1 U11254 ( .A(n10854), .B(n10855), .Y(n11521) );
  inv_1 U11255 ( .A(n11513), .Y(n10855) );
  inv_1 U11256 ( .A(n10854), .Y(n11514) );
  a22oi_1 U11257 ( .A1(n11522), .A2(n11523), .B1(n11524), .B2(n23800), .Y(
        n10854) );
  or2_0 U11258 ( .A(n11523), .B(n11522), .X(n11524) );
  xnor2_1 U11259 ( .A(n11525), .B(n11526), .Y(n11522) );
  xor2_1 U11260 ( .A(n11527), .B(n23769), .X(n11513) );
  nand2_1 U11261 ( .A(n11509), .B(n11511), .Y(n11527) );
  nand2_1 U11262 ( .A(n11528), .B(n10845), .Y(n11511) );
  or2_0 U11263 ( .A(n10845), .B(n11528), .X(n11509) );
  inv_1 U11264 ( .A(n10847), .Y(n10845) );
  nand2_1 U11265 ( .A(inData[30]), .B(n23885), .Y(n11501) );
  o32ai_1 U11266 ( .A1(n11107), .A2(n11529), .A3(n10832), .B1(n11530), .B2(
        n10833), .Y(n10529) );
  xor2_1 U11267 ( .A(n11531), .B(n23687), .X(n11530) );
  xor2_1 U11268 ( .A(n11532), .B(n12452), .X(n11529) );
  or2_0 U11269 ( .A(n10860), .B(n23801), .X(n11532) );
  inv_1 U11270 ( .A(n23885), .Y(n10860) );
  nand2_1 U11271 ( .A(n11533), .B(n11534), .Y(n10528) );
  mux2i_1 U11272 ( .A0(n11535), .A1(n11536), .S(n11537), .Y(n11533) );
  xor2_1 U11273 ( .A(n11538), .B(n11539), .X(n11536) );
  xor2_1 U11274 ( .A(n11540), .B(n11541), .X(n11539) );
  nand2_1 U11275 ( .A(n11542), .B(inData[0]), .Y(n11535) );
  xor2_1 U11276 ( .A(n11543), .B(n11544), .X(n11542) );
  xor2_1 U11277 ( .A(n23971), .B(n23925), .X(n11544) );
  or2_0 U11278 ( .A(n23924), .B(n23706), .X(n11543) );
  o32ai_1 U11279 ( .A1(n11545), .A2(n11546), .A3(n11150), .B1(n11152), .B2(
        n11547), .Y(n10527) );
  xnor2_1 U11280 ( .A(n11548), .B(n11549), .Y(n11547) );
  xor2_1 U11281 ( .A(n23969), .B(n11550), .X(n11549) );
  xor2_1 U11282 ( .A(n11343), .B(n12520), .X(n11546) );
  nand2_1 U11283 ( .A(n23922), .B(n11551), .Y(n10526) );
  xor2_1 U11284 ( .A(n11552), .B(n11553), .X(n11551) );
  xor2_1 U11285 ( .A(n11554), .B(n11555), .X(n11553) );
  nand2_1 U11286 ( .A(n11556), .B(n11557), .Y(n11552) );
  nor2_1 U11287 ( .A(_____9___34419), .B(n11558), .Y(n10525) );
  nand2_1 U11288 ( .A(n11559), .B(n11534), .Y(n10524) );
  mux2i_1 U11289 ( .A0(n11560), .A1(n11561), .S(n11537), .Y(n11559) );
  xnor2_1 U11290 ( .A(n11562), .B(n11563), .Y(n11561) );
  xor2_1 U11291 ( .A(n11564), .B(n11565), .X(n11563) );
  nand2_1 U11292 ( .A(n23925), .B(inData[26]), .Y(n11560) );
  mux4_2 U11293 ( .A0(n11566), .A1(n11567), .A2(n11567), .A3(n11566), .S0(
        n11568), .S1(n11569), .X(n10523) );
  xor2_1 U11294 ( .A(n23706), .B(n11570), .X(n11569) );
  nand2_1 U11295 ( .A(n11571), .B(n23922), .Y(n10522) );
  xor2_1 U11296 ( .A(n11572), .B(n11573), .X(n11571) );
  xor2_1 U11297 ( .A(n11574), .B(n11575), .X(n11573) );
  nand2_1 U11298 ( .A(n11576), .B(n11577), .Y(n11572) );
  xor2_1 U11299 ( .A(n11520), .B(n11578), .X(n11576) );
  or2_0 U11300 ( .A(n47), .B(n11558), .X(n10521) );
  mux2i_1 U11301 ( .A0(n11579), .A1(n11580), .S(n11418), .Y(n10520) );
  a22oi_1 U11302 ( .A1(n11581), .A2(n11582), .B1(n11583), .B2(n11584), .Y(
        n11580) );
  o21ai_0 U11303 ( .A1(n11585), .A2(n11586), .B1(n11584), .Y(n11581) );
  nor3_1 U11304 ( .A(n11587), .B(n10922), .C(n11330), .Y(n11579) );
  xor2_1 U11305 ( .A(n23772), .B(n23681), .X(n11587) );
  nand2_1 U11306 ( .A(n11588), .B(n11503), .Y(n10519) );
  xor2_1 U11307 ( .A(n11589), .B(n11590), .X(n11588) );
  xor2_1 U11308 ( .A(n11591), .B(n55), .X(n11589) );
  nand2_1 U11309 ( .A(n11592), .B(n11593), .Y(n10518) );
  mux2i_1 U11310 ( .A0(n11594), .A1(n11595), .S(n10819), .Y(n11592) );
  xor2_1 U11311 ( .A(n11596), .B(n11597), .X(n11595) );
  xor2_1 U11312 ( .A(n23851), .B(n12579), .X(n11597) );
  nand2_1 U11313 ( .A(n23797), .B(n11598), .Y(n11596) );
  xor2_1 U11314 ( .A(n11599), .B(n11600), .X(n11594) );
  xnor2_1 U11315 ( .A(n23772), .B(n11601), .Y(n11600) );
  xor2_1 U11316 ( .A(n11602), .B(n11603), .X(n11599) );
  nand2_1 U11317 ( .A(n11604), .B(n11500), .Y(n10517) );
  mux2i_1 U11318 ( .A0(n11605), .A1(n11606), .S(n11503), .Y(n11604) );
  xor2_1 U11319 ( .A(n11607), .B(n11608), .X(n11606) );
  xor2_1 U11320 ( .A(n11609), .B(n11610), .X(n11608) );
  xor2_1 U11321 ( .A(n11611), .B(n11612), .X(n11607) );
  nand2_1 U11322 ( .A(n11613), .B(inData[2]), .Y(n11605) );
  xnor2_1 U11323 ( .A(n60), .B(n11614), .Y(n11613) );
  mux2i_1 U11324 ( .A0(n11615), .A1(n11616), .S(n11617), .Y(n10516) );
  a211oi_1 U11325 ( .A1(n23803), .A2(n23804), .B1(n11174), .C1(n11614), .Y(
        n11616) );
  nand2_1 U11326 ( .A(inData[26]), .B(n11618), .Y(n11174) );
  xor2_1 U11327 ( .A(n11619), .B(n11620), .X(n11615) );
  xor2_1 U11328 ( .A(n11621), .B(n11622), .X(n11620) );
  xnor2_1 U11329 ( .A(n11623), .B(n11624), .Y(n11619) );
  nand2_1 U11330 ( .A(n11625), .B(n11626), .Y(n10515) );
  mux2i_1 U11331 ( .A0(n11627), .A1(n11628), .S(n11629), .Y(n11625) );
  xor2_1 U11332 ( .A(n11630), .B(n11631), .X(n11628) );
  xor2_1 U11333 ( .A(n11632), .B(n59), .X(n11630) );
  nand2_1 U11334 ( .A(n11633), .B(n11390), .Y(n10514) );
  mux2i_1 U11335 ( .A0(n11634), .A1(n11635), .S(n11393), .Y(n11633) );
  xor2_1 U11336 ( .A(n11636), .B(n69), .X(n11635) );
  xnor2_1 U11337 ( .A(n11637), .B(n11638), .Y(n11634) );
  o21ai_0 U11338 ( .A1(n11639), .A2(n11640), .B1(n11641), .Y(n11638) );
  mux2i_1 U11339 ( .A0(n11642), .A1(n11643), .S(n11393), .Y(n10513) );
  nand3_1 U11340 ( .A(n11644), .B(n11645), .C(inData[16]), .Y(n11643) );
  xor2_1 U11341 ( .A(n11636), .B(n23937), .X(n11644) );
  xor2_1 U11342 ( .A(n11646), .B(n11647), .X(n11642) );
  mux2i_1 U11343 ( .A0(n11648), .A1(n11649), .S(n11650), .Y(n11647) );
  xnor2_1 U11344 ( .A(n11651), .B(n11652), .Y(n11649) );
  a21oi_1 U11345 ( .A1(n11652), .A2(n11651), .B1(n11653), .Y(n11648) );
  mux2i_1 U11346 ( .A0(n11654), .A1(n11655), .S(n11393), .Y(n10512) );
  o211ai_1 U11347 ( .A1(n70), .A2(n11656), .B1(n11645), .C1(n11636), .Y(n11655) );
  nand2_1 U11348 ( .A(n70), .B(n11656), .Y(n11636) );
  inv_1 U11349 ( .A(n23921), .Y(n11656) );
  xor2_1 U11350 ( .A(n11657), .B(n11658), .X(n11654) );
  xnor2_1 U11351 ( .A(n11659), .B(n11660), .Y(n11658) );
  o22ai_1 U11352 ( .A1(n11661), .A2(n11480), .B1(n11482), .B2(n11662), .Y(
        n10511) );
  xor2_1 U11353 ( .A(n11663), .B(n11664), .X(n11662) );
  xor2_1 U11354 ( .A(n11665), .B(n11666), .X(n11664) );
  xor2_1 U11355 ( .A(n11667), .B(n11668), .X(n11663) );
  nand2_1 U11356 ( .A(n23922), .B(n11669), .Y(n10510) );
  xnor2_1 U11357 ( .A(n10969), .B(n11670), .Y(n11669) );
  xor2_1 U11358 ( .A(n10970), .B(n10968), .X(n11670) );
  inv_1 U11359 ( .A(n11671), .Y(n10968) );
  o21ai_0 U11360 ( .A1(n11672), .A2(n11673), .B1(n11674), .Y(n11671) );
  xor2_1 U11361 ( .A(n11675), .B(n11676), .X(n10969) );
  xor2_1 U11362 ( .A(n11677), .B(n10974), .X(n11676) );
  o22ai_1 U11363 ( .A1(n11678), .A2(n11679), .B1(n11680), .B2(n10629), .Y(
        n10974) );
  and2_0 U11364 ( .A(n11679), .B(n11678), .X(n11680) );
  xor2_1 U11365 ( .A(n10629), .B(n12318), .X(n11675) );
  o22ai_1 U11366 ( .A1(_____90__34411), .A2(n10924), .B1(n11681), .B2(n11420), 
        .Y(n10509) );
  nand2_1 U11367 ( .A(inData[24]), .B(n11495), .Y(n11420) );
  nor2_1 U11368 ( .A(n10774), .B(n11682), .Y(n10508) );
  xor2_1 U11369 ( .A(n11683), .B(n11672), .X(n11682) );
  xor2_1 U11370 ( .A(n11684), .B(n11685), .X(n11672) );
  a21oi_1 U11371 ( .A1(n11490), .A2(n11493), .B1(n11492), .Y(n11685) );
  xor2_1 U11372 ( .A(n11520), .B(n11686), .X(n11492) );
  nor2_1 U11373 ( .A(n11687), .B(n11688), .Y(n11686) );
  nand2_1 U11374 ( .A(n11688), .B(n11687), .Y(n11493) );
  xnor2_1 U11375 ( .A(n11689), .B(n11690), .Y(n11688) );
  xor2_1 U11376 ( .A(n779), .B(n12467), .X(n11690) );
  o21ai_0 U11377 ( .A1(n11691), .A2(n11692), .B1(n11693), .Y(n11490) );
  inv_1 U11378 ( .A(n11694), .Y(n11692) );
  nor2_1 U11379 ( .A(n11695), .B(n11673), .Y(n11683) );
  xor2_1 U11380 ( .A(n11684), .B(n11696), .X(n11673) );
  nor2_1 U11381 ( .A(n11697), .B(n11698), .Y(n11696) );
  inv_1 U11382 ( .A(n11674), .Y(n11695) );
  nand2_1 U11383 ( .A(n11697), .B(n11698), .Y(n11674) );
  xor2_1 U11384 ( .A(n11678), .B(n11699), .X(n11698) );
  xor2_1 U11385 ( .A(n20749), .B(n12467), .X(n11699) );
  a22oi_1 U11386 ( .A1(n11679), .A2(n11689), .B1(n11700), .B2(n779), .Y(n11678) );
  or2_0 U11387 ( .A(n11689), .B(n11679), .X(n11700) );
  o22ai_1 U11388 ( .A1(n12429), .A2(n11701), .B1(n779), .B2(n11702), .Y(n11689) );
  and2_0 U11389 ( .A(n12429), .B(n11701), .X(n11702) );
  o21ai_0 U11390 ( .A1(n11703), .A2(n11498), .B1(n11704), .Y(n10507) );
  nand2_1 U11391 ( .A(__________0_______18822), .B(n11418), .Y(n11704) );
  nor2_1 U11392 ( .A(n10802), .B(n11705), .Y(n10506) );
  xor2_1 U11393 ( .A(n11706), .B(n11707), .X(n11705) );
  xnor2_1 U11394 ( .A(n11708), .B(n11709), .Y(n11707) );
  xor2_1 U11395 ( .A(n11710), .B(n11711), .X(n11706) );
  mux2i_1 U11396 ( .A0(n11712), .A1(n11713), .S(n10819), .Y(n10505) );
  a211oi_1 U11397 ( .A1(n23721), .A2(n11508), .B1(n10821), .C1(n10823), .Y(
        n11713) );
  xor2_1 U11398 ( .A(n11714), .B(n11715), .X(n11712) );
  xnor2_1 U11399 ( .A(n11716), .B(n15), .Y(n11714) );
  nand2_1 U11400 ( .A(n11717), .B(n11500), .Y(n10504) );
  mux2i_1 U11401 ( .A0(n11718), .A1(n11719), .S(n11503), .Y(n11717) );
  xor2_1 U11402 ( .A(n11515), .B(n11720), .X(n11719) );
  xor2_1 U11403 ( .A(n11516), .B(n11519), .X(n11720) );
  a22oi_1 U11404 ( .A1(n11610), .A2(n11609), .B1(n11611), .B2(n11721), .Y(
        n11519) );
  or2_0 U11405 ( .A(n11609), .B(n11610), .X(n11721) );
  or2_0 U11406 ( .A(n11722), .B(n11723), .X(n11611) );
  a21oi_1 U11407 ( .A1(n11724), .A2(n11725), .B1(n12579), .Y(n11723) );
  xor2_1 U11408 ( .A(n11414), .B(n11726), .X(n11722) );
  nor2_1 U11409 ( .A(n11724), .B(n11725), .Y(n11726) );
  inv_1 U11410 ( .A(n11727), .Y(n11724) );
  mux2i_1 U11411 ( .A0(n11728), .A1(n11729), .S(n23799), .Y(n11609) );
  o21ai_0 U11412 ( .A1(n11603), .A2(n11730), .B1(n11731), .Y(n11729) );
  xor2_1 U11413 ( .A(n11603), .B(n11730), .X(n11728) );
  mux2i_1 U11414 ( .A0(n11732), .A1(n11733), .S(n11734), .Y(n11610) );
  nor2_1 U11415 ( .A(n11735), .B(n11736), .Y(n11733) );
  inv_1 U11416 ( .A(n11737), .Y(n11736) );
  o22ai_1 U11417 ( .A1(n11737), .A2(n11738), .B1(n11739), .B2(n11740), .Y(
        n11732) );
  and2_0 U11418 ( .A(n11738), .B(n11737), .X(n11739) );
  o22ai_1 U11419 ( .A1(n11603), .A2(n11730), .B1(n23799), .B2(n11741), .Y(
        n11516) );
  xor2_1 U11420 ( .A(n11742), .B(n11731), .X(n11741) );
  nand2_1 U11421 ( .A(n11603), .B(n11730), .Y(n11731) );
  nand2_1 U11422 ( .A(n11743), .B(n11744), .Y(n11730) );
  xor2_1 U11423 ( .A(n11346), .B(n11745), .X(n11743) );
  nor2_1 U11424 ( .A(n11746), .B(n11747), .Y(n11745) );
  xor2_1 U11425 ( .A(n11748), .B(n11749), .X(n11515) );
  xor2_1 U11426 ( .A(n23800), .B(n12297), .X(n11749) );
  xor2_1 U11427 ( .A(n11523), .B(n11526), .X(n11748) );
  a21oi_1 U11428 ( .A1(outData[31]), .A2(n11750), .B1(n10847), .Y(n11526) );
  nor2_1 U11429 ( .A(n11750), .B(outData[31]), .Y(n10847) );
  inv_1 U11430 ( .A(n11744), .Y(n11750) );
  xor2_1 U11431 ( .A(n11751), .B(n11752), .X(n11744) );
  and2_0 U11432 ( .A(n11746), .B(n11747), .X(n11752) );
  nand2_1 U11433 ( .A(n11753), .B(n10646), .Y(n11718) );
  xnor2_1 U11434 ( .A(n59), .B(n11614), .Y(n11753) );
  nor2_1 U11435 ( .A(n23803), .B(n23804), .Y(n11614) );
  nor2_1 U11436 ( .A(n10774), .B(n11754), .Y(n10503) );
  xor2_1 U11437 ( .A(n11755), .B(n11756), .X(n11754) );
  xor2_1 U11438 ( .A(n11757), .B(n60), .X(n11756) );
  nand2_1 U11439 ( .A(n11758), .B(n11114), .Y(n10502) );
  mux2i_1 U11440 ( .A0(n11759), .A1(n11760), .S(n11117), .Y(n11758) );
  nand2_1 U11441 ( .A(inData[14]), .B(n11761), .Y(n11760) );
  xor2_1 U11442 ( .A(n12476), .B(n11762), .X(n11761) );
  nor2_1 U11443 ( .A(n12522), .B(n818), .Y(n11762) );
  xor2_1 U11444 ( .A(n11763), .B(n11764), .X(n11759) );
  xor2_1 U11445 ( .A(n11765), .B(n23804), .X(n11764) );
  o32ai_1 U11446 ( .A1(n11472), .A2(n10639), .A3(n11330), .B1(n11470), .B2(
        n11766), .Y(n10501) );
  xnor2_1 U11447 ( .A(n11767), .B(n11768), .Y(n11766) );
  a21oi_1 U11448 ( .A1(n11769), .A2(n11770), .B1(n11771), .Y(n11768) );
  mux2i_1 U11449 ( .A0(n11772), .A1(n11773), .S(n11470), .Y(n10500) );
  nor3_1 U11450 ( .A(n11774), .B(n11775), .C(n11472), .Y(n11773) );
  xor2_1 U11451 ( .A(n11776), .B(n11474), .X(n11774) );
  a21oi_1 U11452 ( .A1(n11777), .A2(n11627), .B1(n11778), .Y(n11772) );
  inv_1 U11453 ( .A(n12521), .Y(n11627) );
  inv_1 U11454 ( .A(n11779), .Y(n11777) );
  nor2_1 U11455 ( .A(n11780), .B(n10774), .Y(n10499) );
  xor2_1 U11456 ( .A(n11781), .B(n11782), .X(n11780) );
  nand2_1 U11457 ( .A(n11783), .B(n11784), .Y(n11781) );
  nand4_1 U11458 ( .A(n11785), .B(n11786), .C(n11787), .D(n11788), .Y(n10498)
         );
  nor4_1 U11459 ( .A(n11789), .B(n11790), .C(n11791), .D(n11792), .Y(n11788)
         );
  nand4_1 U11460 ( .A(n11793), .B(n11794), .C(n11795), .D(n11796), .Y(n11789)
         );
  nor4_1 U11461 ( .A(n11797), .B(n11798), .C(n11799), .D(n11800), .Y(n11787)
         );
  and4_1 U11462 ( .A(n11801), .B(n11802), .C(n11803), .D(n11804), .X(n11800)
         );
  and4_1 U11463 ( .A(n11805), .B(n11806), .C(n11807), .D(n11808), .X(n11799)
         );
  a21oi_1 U11464 ( .A1(n11809), .A2(n11810), .B1(n11811), .Y(n11798) );
  o221ai_1 U11465 ( .A1(n11812), .A2(n11813), .B1(n11814), .B2(n11815), .C1(
        n11816), .Y(n11797) );
  o21ai_0 U11466 ( .A1(n11817), .A2(n11818), .B1(n11819), .Y(n11816) );
  and3_1 U11467 ( .A(n11820), .B(n11821), .C(n11822), .X(n11817) );
  nor4_1 U11468 ( .A(n11823), .B(n11824), .C(n11825), .D(n11826), .Y(n11786)
         );
  o221ai_1 U11469 ( .A1(n11827), .A2(n11828), .B1(n11829), .B2(n11830), .C1(
        n11831), .Y(n11823) );
  nor4_1 U11470 ( .A(n11832), .B(n11833), .C(n11834), .D(n11835), .Y(n11785)
         );
  mux2i_1 U11471 ( .A0(n11836), .A1(n11837), .S(n11838), .Y(n11833) );
  and2_0 U11472 ( .A(n11839), .B(n11840), .X(n11837) );
  nor2_1 U11473 ( .A(n11841), .B(n11842), .Y(n11836) );
  o32ai_1 U11474 ( .A1(n11843), .A2(n11844), .A3(n11845), .B1(n11846), .B2(
        n11847), .Y(n11842) );
  or3_1 U11475 ( .A(n11848), .B(n11849), .C(n11850), .X(n11832) );
  inv_1 U11476 ( .A(n11851), .Y(n11849) );
  nand4_1 U11477 ( .A(n11852), .B(n11853), .C(n11854), .D(n11855), .Y(n10497)
         );
  nor4_1 U11478 ( .A(n11856), .B(n11857), .C(n11858), .D(n11859), .Y(n11855)
         );
  inv_1 U11479 ( .A(n11860), .Y(n11859) );
  or3_1 U11480 ( .A(n11861), .B(n11862), .C(n11863), .X(n11857) );
  nand4_1 U11481 ( .A(n11864), .B(n11865), .C(n11866), .D(n11867), .Y(n11856)
         );
  inv_1 U11482 ( .A(n11868), .Y(n11867) );
  a21oi_1 U11483 ( .A1(n11869), .A2(n11870), .B1(n11871), .Y(n11866) );
  nor4_1 U11484 ( .A(n11872), .B(n11873), .C(n11874), .D(n11875), .Y(n11854)
         );
  nand3_1 U11485 ( .A(n11876), .B(n11877), .C(n11878), .Y(n11872) );
  a222oi_1 U11486 ( .A1(n11879), .A2(n11880), .B1(n11881), .B2(n11882), .C1(
        n11838), .C2(n11883), .Y(n11853) );
  a22oi_1 U11487 ( .A1(n11884), .A2(n11885), .B1(n11886), .B2(n11814), .Y(
        n11852) );
  nand3_1 U11488 ( .A(n11887), .B(n11888), .C(n11889), .Y(n10496) );
  nor4_1 U11489 ( .A(n11890), .B(n11891), .C(n11892), .D(n11893), .Y(n11889)
         );
  nand3_1 U11490 ( .A(n11796), .B(n11894), .C(n11895), .Y(n11891) );
  inv_1 U11491 ( .A(n11896), .Y(n11796) );
  a21oi_1 U11492 ( .A1(n11897), .A2(n11898), .B1(n11838), .Y(n11896) );
  o221ai_1 U11493 ( .A1(n11805), .A2(n11899), .B1(n11900), .B2(n11901), .C1(
        n11902), .Y(n11890) );
  a222oi_1 U11494 ( .A1(n11790), .A2(n11870), .B1(n11903), .B2(n11827), .C1(
        n11904), .C2(n11905), .Y(n11902) );
  nor3_1 U11495 ( .A(n11906), .B(n11907), .C(n11908), .Y(n11888) );
  nand3_1 U11496 ( .A(n11909), .B(n11910), .C(n11864), .Y(n11906) );
  a21oi_1 U11497 ( .A1(n11819), .A2(n11911), .B1(n11912), .Y(n11864) );
  nor4_1 U11498 ( .A(n11913), .B(n11914), .C(n11915), .D(n11916), .Y(n11887)
         );
  or3_1 U11499 ( .A(n11917), .B(n11918), .C(n11919), .X(n10495) );
  nand4_1 U11500 ( .A(n11920), .B(n11921), .C(n11922), .D(n11923), .Y(n11919)
         );
  nor4_1 U11501 ( .A(n11924), .B(n11925), .C(n11926), .D(n11927), .Y(n11923)
         );
  o22ai_1 U11502 ( .A1(n11829), .A2(n11928), .B1(n11819), .B2(n11929), .Y(
        n11925) );
  nor3_1 U11503 ( .A(n11930), .B(n11931), .C(n11932), .Y(n11922) );
  inv_1 U11504 ( .A(n11933), .Y(n11921) );
  inv_1 U11505 ( .A(n11934), .Y(n11920) );
  o221ai_1 U11506 ( .A1(n11935), .A2(n11870), .B1(n11905), .B2(n11936), .C1(
        n11937), .Y(n11918) );
  a222oi_1 U11507 ( .A1(n11938), .A2(n11884), .B1(n11939), .B2(n11900), .C1(
        n11940), .C2(n11827), .Y(n11937) );
  inv_1 U11508 ( .A(n11846), .Y(n11939) );
  inv_1 U11509 ( .A(n11941), .Y(n11938) );
  nand4_1 U11510 ( .A(n11840), .B(n11942), .C(n11943), .D(n11944), .Y(n11917)
         );
  nor3_1 U11511 ( .A(n11945), .B(n11892), .C(n11792), .Y(n11944) );
  inv_1 U11512 ( .A(n11830), .Y(n11892) );
  nand4_1 U11513 ( .A(n11946), .B(n11947), .C(n11948), .D(n11949), .Y(n10494)
         );
  nor3_1 U11514 ( .A(n11950), .B(n11940), .C(n11951), .Y(n11949) );
  a21oi_1 U11515 ( .A1(n11952), .A2(n11943), .B1(n11953), .Y(n11951) );
  nand3_1 U11516 ( .A(n11954), .B(n11955), .C(n11956), .Y(n11950) );
  a221oi_1 U11517 ( .A1(n11957), .A2(n11958), .B1(n11959), .B2(n11882), .C1(
        n11960), .Y(n11948) );
  o22ai_1 U11518 ( .A1(n11900), .A2(n11876), .B1(n11905), .B2(n11961), .Y(
        n11960) );
  nor4_1 U11519 ( .A(n11862), .B(n11962), .C(n11963), .D(n11914), .Y(n11947)
         );
  o221ai_1 U11520 ( .A1(n11905), .A2(n11964), .B1(n11819), .B2(n11965), .C1(
        n11966), .Y(n11914) );
  a211oi_1 U11521 ( .A1(n11967), .A2(n11884), .B1(n11968), .C1(n11969), .Y(
        n11966) );
  o21ai_0 U11522 ( .A1(n11819), .A2(n11970), .B1(n11851), .Y(n11962) );
  a221oi_1 U11523 ( .A1(n11814), .A2(n11971), .B1(n11953), .B2(n11972), .C1(
        n11973), .Y(n11851) );
  o21ai_0 U11524 ( .A1(n11974), .A2(n11811), .B1(n11975), .Y(n11973) );
  nand4_1 U11525 ( .A(n11909), .B(n11976), .C(n11977), .D(n11978), .Y(n11862)
         );
  nor4_1 U11526 ( .A(n11979), .B(n11980), .C(n11981), .D(n11982), .Y(n11978)
         );
  inv_1 U11527 ( .A(n11983), .Y(n11981) );
  nand3_1 U11528 ( .A(n11984), .B(n11898), .C(n11985), .Y(n11979) );
  a221oi_1 U11529 ( .A1(n11986), .A2(n11900), .B1(n11987), .B2(n11988), .C1(
        n11989), .Y(n11977) );
  a21oi_1 U11530 ( .A1(n11990), .A2(n11991), .B1(n11805), .Y(n11989) );
  inv_1 U11531 ( .A(n11992), .Y(n11976) );
  a211oi_1 U11532 ( .A1(n11993), .A2(n11838), .B1(n11994), .C1(n11945), .Y(
        n11909) );
  nor4_1 U11533 ( .A(n11995), .B(n11996), .C(n11997), .D(n11998), .Y(n11946)
         );
  mux2i_1 U11534 ( .A0(n11999), .A1(n11813), .S(n11812), .Y(n11998) );
  nor2_1 U11535 ( .A(n12000), .B(n12001), .Y(n11813) );
  inv_1 U11536 ( .A(n12002), .Y(n12001) );
  nor3_1 U11537 ( .A(n12003), .B(n12004), .C(n11893), .Y(n11999) );
  inv_1 U11538 ( .A(n12005), .Y(n11996) );
  nand3_1 U11539 ( .A(n12006), .B(n12007), .C(n12008), .Y(n10493) );
  nor4_1 U11540 ( .A(n12009), .B(n12010), .C(n12011), .D(n12012), .Y(n12008)
         );
  inv_1 U11541 ( .A(n11928), .Y(n12012) );
  nand3_1 U11542 ( .A(n11941), .B(n12013), .C(n11970), .Y(n12010) );
  nand3_1 U11543 ( .A(n11983), .B(n12014), .C(n12015), .Y(n12009) );
  a21oi_1 U11544 ( .A1(n12016), .A2(n11953), .B1(n12017), .Y(n12015) );
  a21oi_1 U11545 ( .A1(n12018), .A2(n12019), .B1(n11905), .Y(n12017) );
  nor4_1 U11546 ( .A(n11912), .B(n12020), .C(n11913), .D(n11931), .Y(n12007)
         );
  nand4_1 U11547 ( .A(n12021), .B(n12022), .C(n12023), .D(n12024), .Y(n11931)
         );
  a211oi_1 U11548 ( .A1(n11986), .A2(n11838), .B1(n12025), .C1(n12026), .Y(
        n12024) );
  a21oi_1 U11549 ( .A1(n12027), .A2(n12028), .B1(n11819), .Y(n12026) );
  inv_1 U11550 ( .A(n12029), .Y(n12023) );
  nand2_1 U11551 ( .A(n11971), .B(n11814), .Y(n12022) );
  inv_1 U11552 ( .A(n12030), .Y(n12021) );
  o22ai_1 U11553 ( .A1(n11880), .A2(n12031), .B1(n11953), .B2(n12032), .Y(
        n11913) );
  o21ai_0 U11554 ( .A1(n11900), .A2(n12033), .B1(n12034), .Y(n12020) );
  inv_1 U11555 ( .A(n11824), .Y(n12034) );
  o221ai_1 U11556 ( .A1(n11953), .A2(n11985), .B1(n11905), .B2(n11984), .C1(
        n11936), .Y(n11824) );
  o211ai_1 U11557 ( .A1(n11953), .A2(n12035), .B1(n12036), .C1(n12037), .Y(
        n11912) );
  nor4_1 U11558 ( .A(n12038), .B(n12039), .C(n12040), .D(n12041), .Y(n12006)
         );
  nand3_1 U11559 ( .A(n12042), .B(n12043), .C(n12044), .Y(n10492) );
  nor4_1 U11560 ( .A(n12045), .B(n12046), .C(n12047), .D(n11972), .Y(n12044)
         );
  inv_1 U11561 ( .A(n12048), .Y(n11972) );
  nand3_1 U11562 ( .A(n11901), .B(n11894), .C(n12031), .Y(n12046) );
  o221ai_1 U11563 ( .A1(n11953), .A2(n11943), .B1(n11814), .B2(n12018), .C1(
        n12049), .Y(n12045) );
  a21oi_1 U11564 ( .A1(n12050), .A2(n11988), .B1(n12051), .Y(n12049) );
  nor4_1 U11565 ( .A(n12052), .B(n11826), .C(n11863), .D(n11930), .Y(n12043)
         );
  o211ai_1 U11566 ( .A1(n11819), .A2(n11965), .B1(n12053), .C1(n12054), .Y(
        n11930) );
  a211oi_1 U11567 ( .A1(n11791), .A2(n11805), .B1(n12055), .C1(n11967), .Y(
        n12054) );
  inv_1 U11568 ( .A(n12056), .Y(n11967) );
  inv_1 U11569 ( .A(n11954), .Y(n12055) );
  or3_1 U11570 ( .A(n12057), .B(n12058), .C(n12059), .X(n11863) );
  o22ai_1 U11571 ( .A1(n12014), .A2(n11827), .B1(n11928), .B2(n11829), .Y(
        n12059) );
  o22ai_1 U11572 ( .A1(n11805), .A2(n11991), .B1(n11880), .B2(n12060), .Y(
        n11826) );
  nor2_1 U11573 ( .A(n11884), .B(n12061), .Y(n12052) );
  nor4_1 U11574 ( .A(n12040), .B(n12062), .C(n12063), .D(n12064), .Y(n12042)
         );
  or4_1 U11575 ( .A(n12065), .B(n11932), .C(n12066), .D(n12067), .X(n12040) );
  or4_1 U11576 ( .A(n12068), .B(n11980), .C(n12069), .D(n11886), .X(n12067) );
  o22ai_1 U11577 ( .A1(n11814), .A2(n12070), .B1(n12071), .B2(n11870), .Y(
        n12068) );
  nor2_1 U11578 ( .A(n12003), .B(n12072), .Y(n12071) );
  o21ai_0 U11579 ( .A1(n11898), .A2(n11838), .B1(n12073), .Y(n12066) );
  nand4_1 U11580 ( .A(n12074), .B(n12075), .C(n12076), .D(n12077), .Y(n11932)
         );
  a221oi_1 U11581 ( .A1(n12078), .A2(n11805), .B1(n12079), .B2(n11838), .C1(
        n12080), .Y(n12077) );
  nand2_1 U11582 ( .A(n11873), .B(n11814), .Y(n12075) );
  inv_1 U11583 ( .A(n11861), .Y(n12074) );
  o22ai_1 U11584 ( .A1(n11953), .A2(n12081), .B1(n11988), .B2(n12082), .Y(
        n11861) );
  a21oi_1 U11585 ( .A1(n12083), .A2(n12084), .B1(n11968), .Y(n12082) );
  nand4_1 U11586 ( .A(n12085), .B(n12086), .C(n12087), .D(n12088), .Y(n10491)
         );
  nor4_1 U11587 ( .A(n12089), .B(n12090), .C(n11848), .D(n11871), .Y(n12088)
         );
  o21ai_0 U11588 ( .A1(n11812), .A2(n12091), .B1(n12092), .Y(n11871) );
  nand4_1 U11589 ( .A(n12093), .B(n12094), .C(n12095), .D(n12096), .Y(n11848)
         );
  and4_1 U11590 ( .A(n12097), .B(n11965), .C(n12098), .D(n12013), .X(n12096)
         );
  inv_1 U11591 ( .A(n12099), .Y(n12097) );
  o32ai_1 U11592 ( .A1(n12100), .A2(n12101), .A3(n11870), .B1(n11811), .B2(
        n12102), .Y(n12099) );
  a22oi_1 U11593 ( .A1(n11911), .A2(n11819), .B1(n11880), .B2(n11994), .Y(
        n12095) );
  inv_1 U11594 ( .A(n12103), .Y(n11994) );
  inv_1 U11595 ( .A(n11956), .Y(n11911) );
  o22ai_1 U11596 ( .A1(n11827), .A2(n11952), .B1(n11805), .B2(n12056), .Y(
        n12090) );
  nand4_1 U11597 ( .A(n12104), .B(n12105), .C(n12106), .D(n11985), .Y(n12089)
         );
  o21ai_0 U11598 ( .A1(n11987), .A2(n12107), .B1(n11819), .Y(n12105) );
  nand2_1 U11599 ( .A(n11812), .B(n11825), .Y(n12104) );
  o21ai_0 U11600 ( .A1(n12108), .A2(n12100), .B1(n12109), .Y(n11825) );
  inv_1 U11601 ( .A(n11807), .Y(n12108) );
  nor4_1 U11602 ( .A(n11908), .B(n11933), .C(n12041), .D(n12110), .Y(n12087)
         );
  nand3_1 U11603 ( .A(n12111), .B(n12112), .C(n12113), .Y(n12041) );
  a21oi_1 U11604 ( .A1(n11790), .A2(n11870), .B1(n12114), .Y(n12113) );
  a21oi_1 U11605 ( .A1(n12048), .A2(n11878), .B1(n11953), .Y(n12114) );
  o221ai_1 U11606 ( .A1(n11882), .A2(n11809), .B1(n11814), .B2(n11964), .C1(
        n12115), .Y(n11933) );
  a21oi_1 U11607 ( .A1(n12116), .A2(n11900), .B1(n11992), .Y(n12115) );
  o22ai_1 U11608 ( .A1(n12117), .A2(n11870), .B1(n11829), .B2(n12060), .Y(
        n11992) );
  o22ai_1 U11609 ( .A1(n11814), .A2(n11984), .B1(n11954), .B2(n11953), .Y(
        n11908) );
  nor2_1 U11610 ( .A(n12118), .B(n12119), .Y(n12085) );
  nand3_1 U11611 ( .A(n12120), .B(n12121), .C(n12122), .Y(n10490) );
  nor4_1 U11612 ( .A(n12123), .B(n12124), .C(n12058), .D(n12125), .Y(n12122)
         );
  nand3_1 U11613 ( .A(n12060), .B(n12126), .C(n12127), .Y(n12124) );
  nand3_1 U11614 ( .A(n12128), .B(n12129), .C(n12130), .Y(n12060) );
  nand4_1 U11615 ( .A(n11810), .B(n11941), .C(n11964), .D(n12131), .Y(n12123)
         );
  a21oi_1 U11616 ( .A1(n12132), .A2(n11905), .B1(n11940), .Y(n12131) );
  inv_1 U11617 ( .A(n12014), .Y(n11940) );
  nor4_1 U11618 ( .A(n12133), .B(n12134), .C(n11850), .D(n11915), .Y(n12121)
         );
  nand4_1 U11619 ( .A(n12135), .B(n12136), .C(n12137), .D(n12138), .Y(n11915)
         );
  and4_1 U11620 ( .A(n12139), .B(n11991), .C(n12140), .D(n12141), .X(n12138)
         );
  and4_1 U11621 ( .A(n11793), .B(n12098), .C(n12142), .D(n11809), .X(n12139)
         );
  nor4_1 U11622 ( .A(n12143), .B(n11980), .C(n12144), .D(n12145), .Y(n12137)
         );
  nor2_1 U11623 ( .A(n11963), .B(n12146), .Y(n12135) );
  o22ai_1 U11624 ( .A1(n11905), .A2(n11936), .B1(n11829), .B2(n12147), .Y(
        n11963) );
  nand3_1 U11625 ( .A(n12148), .B(n12149), .C(n12150), .Y(n11850) );
  nor4_1 U11626 ( .A(n12151), .B(n12152), .C(n11904), .D(n11875), .Y(n12150)
         );
  a22oi_1 U11627 ( .A1(n12047), .A2(n11988), .B1(n11812), .B2(n12153), .Y(
        n12148) );
  inv_1 U11628 ( .A(n12154), .Y(n12153) );
  o21ai_0 U11629 ( .A1(n11812), .A2(n11935), .B1(n12155), .Y(n12134) );
  inv_1 U11630 ( .A(n12094), .Y(n12133) );
  nor3_1 U11631 ( .A(n12004), .B(n12050), .C(n11903), .Y(n12094) );
  inv_1 U11632 ( .A(n12156), .Y(n11903) );
  nor4_1 U11633 ( .A(n12157), .B(n12158), .C(n11995), .D(n12118), .Y(n12120)
         );
  nand4_1 U11634 ( .A(n12036), .B(n11974), .C(n12159), .D(n12160), .Y(n12118)
         );
  a222oi_1 U11635 ( .A1(n12161), .A2(n11827), .B1(n12079), .B2(n11900), .C1(
        n12162), .C2(n11884), .Y(n12160) );
  inv_1 U11636 ( .A(n11876), .Y(n12079) );
  nor2_1 U11637 ( .A(n12163), .B(n10730), .Y(n12159) );
  nand2_1 U11638 ( .A(n12164), .B(n12165), .Y(n12157) );
  mux2i_1 U11639 ( .A0(n12166), .A1(n12167), .S(n11827), .Y(n12165) );
  nand2_1 U11640 ( .A(n12037), .B(n12032), .Y(n12166) );
  mux2i_1 U11641 ( .A0(n12080), .A1(n11969), .S(n11884), .Y(n12164) );
  nand3_1 U11642 ( .A(n12168), .B(n12169), .C(n12170), .Y(n10489) );
  nor4_1 U11643 ( .A(n12171), .B(n12172), .C(n12173), .D(n12174), .Y(n12170)
         );
  a21oi_1 U11644 ( .A1(n12014), .A2(n12035), .B1(n11827), .Y(n12174) );
  a21oi_1 U11645 ( .A1(n11846), .A2(n11897), .B1(n11900), .Y(n12173) );
  o22ai_1 U11646 ( .A1(n12175), .A2(n11884), .B1(n11814), .B2(n11865), .Y(
        n12172) );
  nor2_1 U11647 ( .A(n11971), .B(n12176), .Y(n11865) );
  nand3_1 U11648 ( .A(n12147), .B(n11970), .C(n12177), .Y(n12171) );
  and3_1 U11649 ( .A(n11984), .B(n12178), .C(n12126), .X(n12177) );
  nor4_1 U11650 ( .A(n11834), .B(n12179), .C(n11835), .D(n12146), .Y(n12169)
         );
  o221ai_1 U11651 ( .A1(n12180), .A2(n11870), .B1(n11827), .B2(n12081), .C1(
        n12102), .Y(n12146) );
  nor2_1 U11652 ( .A(n11792), .B(n12003), .Y(n12180) );
  inv_1 U11653 ( .A(n12181), .Y(n11792) );
  nand4_1 U11654 ( .A(n11895), .B(n12182), .C(n12183), .D(n12184), .Y(n11835)
         );
  a211oi_1 U11655 ( .A1(n11827), .A2(n12185), .B1(n11924), .C1(n12186), .Y(
        n12184) );
  inv_1 U11656 ( .A(n12155), .Y(n12186) );
  a221oi_1 U11657 ( .A1(n11874), .A2(n11884), .B1(n11945), .B2(n11814), .C1(
        n12187), .Y(n12155) );
  o21ai_0 U11658 ( .A1(n11954), .A2(n11827), .B1(n12188), .Y(n12187) );
  inv_1 U11659 ( .A(n12189), .Y(n11945) );
  o211ai_1 U11660 ( .A1(n11884), .A2(n12190), .B1(n12019), .C1(n12191), .Y(
        n11924) );
  inv_1 U11661 ( .A(n12192), .Y(n12185) );
  o22ai_1 U11662 ( .A1(n11988), .A2(n11965), .B1(n11870), .B2(n12193), .Y(
        n12179) );
  nand4_1 U11663 ( .A(n12140), .B(n11955), .C(n12027), .D(n12194), .Y(n11834)
         );
  nor3_1 U11664 ( .A(n12195), .B(n11879), .C(n12196), .Y(n12194) );
  a21oi_1 U11665 ( .A1(n11901), .A2(n12141), .B1(n11900), .Y(n12196) );
  inv_1 U11666 ( .A(n12031), .Y(n11879) );
  a21oi_1 U11667 ( .A1(n11990), .A2(n12197), .B1(n11805), .Y(n12195) );
  inv_1 U11668 ( .A(n12163), .Y(n11955) );
  nor2_1 U11669 ( .A(n12033), .B(n11838), .Y(n12163) );
  nor4_1 U11670 ( .A(n11916), .B(n12029), .C(n11997), .D(n12119), .Y(n12168)
         );
  nand4_1 U11671 ( .A(n12198), .B(n12005), .C(n12199), .D(n12200), .Y(n12119)
         );
  nor3_1 U11672 ( .A(n12201), .B(n11881), .C(n12016), .Y(n12200) );
  o21ai_0 U11673 ( .A1(n11953), .A2(n12032), .B1(n12202), .Y(n12201) );
  a21oi_1 U11674 ( .A1(n11838), .A2(n12203), .B1(n12204), .Y(n12199) );
  nor3_1 U11675 ( .A(n12152), .B(n12011), .C(n12205), .Y(n12005) );
  o22ai_1 U11676 ( .A1(n11805), .A2(n11899), .B1(n11880), .B2(n12206), .Y(
        n12205) );
  and3_1 U11677 ( .A(n11988), .B(n12084), .C(n12083), .X(n12152) );
  nand4_1 U11678 ( .A(n12127), .B(n12013), .C(n12156), .D(n12207), .Y(n11997)
         );
  a22oi_1 U11679 ( .A1(n12050), .A2(n11819), .B1(n12162), .B2(n11805), .Y(
        n12207) );
  and2_0 U11680 ( .A(n12083), .B(n12208), .X(n12050) );
  and2_0 U11681 ( .A(n12209), .B(n11958), .X(n12083) );
  nand2_1 U11682 ( .A(n11869), .B(n11812), .Y(n12013) );
  inv_1 U11683 ( .A(n12025), .Y(n12127) );
  nor2_1 U11684 ( .A(n12091), .B(n11870), .Y(n12025) );
  o22ai_1 U11685 ( .A1(n11905), .A2(n11961), .B1(n11819), .B2(n11956), .Y(
        n12029) );
  nand4_1 U11686 ( .A(n12112), .B(n11975), .C(n12210), .D(n12211), .Y(n11916)
         );
  a221oi_1 U11687 ( .A1(n12151), .A2(n11884), .B1(n11982), .B2(n11988), .C1(
        n12167), .Y(n12211) );
  inv_1 U11688 ( .A(n12061), .Y(n12151) );
  a21oi_1 U11689 ( .A1(n12069), .A2(n11811), .B1(n12004), .Y(n12210) );
  inv_1 U11690 ( .A(n12212), .Y(n12004) );
  nand4_1 U11691 ( .A(n12213), .B(n12214), .C(n12215), .D(n12216), .Y(n10488)
         );
  nor4_1 U11692 ( .A(n12217), .B(n12038), .C(n11926), .D(n12065), .Y(n12216)
         );
  o221ai_1 U11693 ( .A1(n12218), .A2(n11900), .B1(n11814), .B2(n12189), .C1(
        n12178), .Y(n12065) );
  nor2_1 U11694 ( .A(n12116), .B(n11993), .Y(n12218) );
  nand2_1 U11695 ( .A(n11839), .B(n12219), .Y(n11993) );
  nand4_1 U11696 ( .A(n12220), .B(n12221), .C(n12222), .D(n12223), .Y(n11839)
         );
  o22ai_1 U11697 ( .A1(n12103), .A2(n11829), .B1(n11900), .B2(n11897), .Y(
        n11926) );
  o21ai_0 U11698 ( .A1(n11884), .A2(n11991), .B1(n12202), .Y(n12038) );
  inv_1 U11699 ( .A(n12144), .Y(n12202) );
  nor2_1 U11700 ( .A(n11840), .B(n11838), .Y(n12144) );
  nand3_1 U11701 ( .A(n12224), .B(n12225), .C(n12226), .Y(n12217) );
  a21oi_1 U11702 ( .A1(n11982), .A2(n11819), .B1(n12227), .Y(n12226) );
  a21oi_1 U11703 ( .A1(n12109), .A2(n12154), .B1(n11870), .Y(n12227) );
  o21ai_0 U11704 ( .A1(n11881), .A2(n12069), .B1(n11811), .Y(n12225) );
  inv_1 U11705 ( .A(n11810), .Y(n11881) );
  o21ai_0 U11706 ( .A1(n12228), .A2(n11873), .B1(n11814), .Y(n12224) );
  nor3_1 U11707 ( .A(n12229), .B(n12230), .C(n12231), .Y(n12215) );
  mux2i_1 U11708 ( .A0(n11990), .A1(n11877), .S(n11884), .Y(n12231) );
  mux2i_1 U11709 ( .A0(n11953), .A1(n12232), .S(n12233), .Y(n12229) );
  nor4_1 U11710 ( .A(n12234), .B(n12235), .C(n12236), .D(n12161), .Y(n12233)
         );
  nand2_1 U11711 ( .A(n11954), .B(n12192), .Y(n12235) );
  nand4_1 U11712 ( .A(n12237), .B(n12037), .C(n11985), .D(n12156), .Y(n12234)
         );
  nand4_1 U11713 ( .A(n12238), .B(n12084), .C(n12239), .D(n11801), .Y(n12156)
         );
  nand4_1 U11714 ( .A(n11840), .B(n11941), .C(n12193), .D(n12240), .Y(n12232)
         );
  nand4_1 U11715 ( .A(n12241), .B(n12242), .C(n12243), .D(n12244), .Y(n12240)
         );
  nor4_1 U11716 ( .A(n12245), .B(n12246), .C(n11791), .D(n11969), .Y(n12244)
         );
  inv_1 U11717 ( .A(n12190), .Y(n11969) );
  nand3_1 U11718 ( .A(n12098), .B(n12142), .C(n11830), .Y(n12246) );
  nand4_1 U11719 ( .A(n12048), .B(n12212), .C(n12247), .D(n12102), .Y(n12245)
         );
  nor2_1 U11720 ( .A(n12057), .B(n12248), .Y(n12247) );
  nor3_1 U11721 ( .A(n12249), .B(n12250), .C(n12162), .Y(n12243) );
  nand3_1 U11722 ( .A(n11936), .B(n11898), .C(n12106), .Y(n12249) );
  nor3_1 U11723 ( .A(n12251), .B(n11885), .C(n11858), .Y(n12242) );
  nor2_1 U11724 ( .A(n12252), .B(n11883), .Y(n12241) );
  inv_1 U11725 ( .A(n12253), .Y(n12214) );
  nor2_1 U11726 ( .A(n12062), .B(n12254), .Y(n12213) );
  nand4_1 U11727 ( .A(n12255), .B(n12256), .C(n12257), .D(n12258), .Y(n12062)
         );
  a221oi_1 U11728 ( .A1(n12143), .A2(n11953), .B1(n12259), .B2(n11882), .C1(
        n12260), .Y(n12258) );
  inv_1 U11729 ( .A(n11907), .Y(n12255) );
  o21ai_0 U11730 ( .A1(n11884), .A2(n11941), .B1(n12183), .Y(n11907) );
  nand4_1 U11731 ( .A(n12261), .B(n12262), .C(n12263), .D(n12264), .Y(n10487)
         );
  and4_1 U11732 ( .A(n12265), .B(n12112), .C(n12098), .D(n12266), .X(n12264)
         );
  nand3_1 U11733 ( .A(n12267), .B(n11821), .C(n12268), .Y(n12098) );
  nand2_1 U11734 ( .A(n12047), .B(n11819), .Y(n12112) );
  and2_0 U11735 ( .A(n12269), .B(n12270), .X(n12047) );
  a21oi_1 U11736 ( .A1(n11819), .A2(n11968), .B1(n11875), .Y(n12265) );
  inv_1 U11737 ( .A(n12206), .Y(n11875) );
  inv_1 U11738 ( .A(n12271), .Y(n11968) );
  a211oi_1 U11739 ( .A1(n12003), .A2(n11870), .B1(n12272), .C1(n12273), .Y(
        n12263) );
  inv_1 U11740 ( .A(n11831), .Y(n12273) );
  a21oi_1 U11741 ( .A1(n11812), .A2(n11893), .B1(n11885), .Y(n11831) );
  o22ai_1 U11742 ( .A1(n11910), .A2(n11900), .B1(n11905), .B2(n11815), .Y(
        n12272) );
  inv_1 U11743 ( .A(n12106), .Y(n12003) );
  nor4_1 U11744 ( .A(n11934), .B(n12039), .C(n12063), .D(n12110), .Y(n12262)
         );
  nand2_1 U11745 ( .A(n11897), .B(n12140), .Y(n12110) );
  nand2_1 U11746 ( .A(n12057), .B(n11819), .Y(n12140) );
  inv_1 U11747 ( .A(n12028), .Y(n12057) );
  nand3_1 U11748 ( .A(n12084), .B(n12274), .C(n12209), .Y(n12028) );
  nand3_1 U11749 ( .A(n12275), .B(n11802), .C(n12276), .Y(n11897) );
  nand4_1 U11750 ( .A(n11810), .B(n12190), .C(n12277), .D(n12278), .Y(n12063)
         );
  a221oi_1 U11751 ( .A1(n11884), .A2(n11874), .B1(n11904), .B2(n11905), .C1(
        n11868), .Y(n12278) );
  o21ai_0 U11752 ( .A1(n11870), .A2(n12212), .B1(n12188), .Y(n11868) );
  nand2_1 U11753 ( .A(n12279), .B(n12280), .Y(n12188) );
  nand3_1 U11754 ( .A(n12128), .B(n12129), .C(n12208), .Y(n12212) );
  inv_1 U11755 ( .A(n11961), .Y(n11904) );
  inv_1 U11756 ( .A(n12281), .Y(n11874) );
  a21oi_1 U11757 ( .A1(n11959), .A2(n11811), .B1(n12282), .Y(n12277) );
  inv_1 U11758 ( .A(n12032), .Y(n12282) );
  nand3_1 U11759 ( .A(n12283), .B(n12084), .C(n12284), .Y(n12032) );
  inv_1 U11760 ( .A(n12102), .Y(n11959) );
  nand3_1 U11761 ( .A(n12270), .B(n12285), .C(n12286), .Y(n12102) );
  nand4_1 U11762 ( .A(n12238), .B(n12208), .C(n11958), .D(n11801), .Y(n11810)
         );
  o22ai_1 U11763 ( .A1(n11812), .A2(n12154), .B1(n11827), .B2(n11954), .Y(
        n12039) );
  nand3_1 U11764 ( .A(n12287), .B(n12288), .C(n12267), .Y(n11954) );
  nand4_1 U11765 ( .A(n11952), .B(n12073), .C(n12289), .D(n12290), .Y(n11934)
         );
  nor4_1 U11766 ( .A(n12291), .B(n12143), .C(n12292), .D(n12260), .Y(n12290)
         );
  inv_1 U11767 ( .A(n12183), .Y(n12292) );
  nand3_1 U11768 ( .A(n11958), .B(n11953), .C(n11957), .Y(n12183) );
  inv_1 U11769 ( .A(n11878), .Y(n12143) );
  o21ai_0 U11770 ( .A1(n11827), .A2(n12293), .B1(n12036), .Y(n12291) );
  nand3_1 U11771 ( .A(n12294), .B(n12221), .C(n12295), .Y(n12036) );
  and3_1 U11772 ( .A(n11814), .B(n12384), .C(n11802), .X(n12295) );
  inv_1 U11773 ( .A(n12167), .Y(n12293) );
  nand2_1 U11774 ( .A(n12048), .B(n11985), .Y(n12167) );
  a21oi_1 U11775 ( .A1(n12069), .A2(n11882), .B1(n12204), .Y(n12289) );
  o21ai_0 U11776 ( .A1(n11953), .A2(n12237), .B1(n11991), .Y(n12204) );
  nand3_1 U11777 ( .A(n12296), .B(n12276), .C(n12298), .Y(n11991) );
  nand4_1 U11778 ( .A(n12221), .B(n12300), .C(n12301), .D(n12384), .Y(n12237)
         );
  inv_1 U11779 ( .A(n11974), .Y(n12069) );
  inv_1 U11780 ( .A(n11995), .Y(n12073) );
  nand2_1 U11781 ( .A(n12197), .B(n12182), .Y(n11995) );
  nand4_1 U11782 ( .A(n12274), .B(n11820), .C(n11882), .D(n11806), .Y(n12182)
         );
  inv_1 U11783 ( .A(n11811), .Y(n11882) );
  nand3_1 U11784 ( .A(inData[30]), .B(n12303), .C(inData[9]), .Y(n11811) );
  inv_1 U11785 ( .A(n12251), .Y(n11952) );
  nor4_1 U11786 ( .A(n11883), .B(n12158), .C(n12230), .D(n12304), .Y(n12261)
         );
  nand4_1 U11787 ( .A(n12136), .B(n12092), .C(n12053), .D(n12306), .Y(n12230)
         );
  a221oi_1 U11788 ( .A1(n11886), .A2(n11905), .B1(n11987), .B2(n11819), .C1(
        n12011), .Y(n12306) );
  inv_1 U11789 ( .A(n12307), .Y(n12011) );
  inv_1 U11790 ( .A(n12027), .Y(n11987) );
  and2_0 U11791 ( .A(n11975), .B(n12309), .X(n12053) );
  nand3_1 U11792 ( .A(n12311), .B(n11808), .C(n12312), .Y(n11975) );
  and3_1 U11793 ( .A(n11988), .B(n11801), .C(n12275), .X(n12312) );
  inv_1 U11794 ( .A(n12313), .Y(n12092) );
  o22ai_1 U11795 ( .A1(n11900), .A2(n11846), .B1(n11880), .B2(n12147), .Y(
        n12313) );
  nand2_1 U11796 ( .A(n12314), .B(n11801), .Y(n12147) );
  nand3_1 U11797 ( .A(n12315), .B(n12317), .C(n11808), .Y(n11846) );
  a22oi_1 U11798 ( .A1(n11870), .A2(n11869), .B1(n11953), .B2(n12016), .Y(
        n12136) );
  inv_1 U11799 ( .A(n11943), .Y(n12016) );
  nand3_1 U11800 ( .A(n11958), .B(n12288), .C(n12287), .Y(n11943) );
  mux2i_1 U11801 ( .A0(n12031), .A1(n12103), .S(n11829), .Y(n12158) );
  nand3_1 U11802 ( .A(n12208), .B(n12128), .C(n12285), .Y(n12031) );
  nand3_1 U11803 ( .A(n11901), .B(n12321), .C(n11840), .Y(n11883) );
  nand3_1 U11804 ( .A(n11822), .B(n12322), .C(n12323), .Y(n11840) );
  nand3_1 U11805 ( .A(n12324), .B(n12325), .C(n12326), .Y(n10486) );
  nor4_1 U11806 ( .A(n12327), .B(n12328), .C(n11886), .D(n11980), .Y(n12326)
         );
  nor4_1 U11807 ( .A(n11843), .B(n11845), .C(n11900), .D(n11844), .Y(n11980)
         );
  inv_1 U11808 ( .A(n12268), .Y(n11845) );
  inv_1 U11809 ( .A(n11964), .Y(n11886) );
  nand3_1 U11810 ( .A(n12315), .B(n12329), .C(n12332), .Y(n11964) );
  nor3_1 U11811 ( .A(n12334), .B(n12335), .C(n11801), .Y(n12332) );
  o22ai_1 U11812 ( .A1(n12175), .A2(n11884), .B1(n12018), .B2(n11905), .Y(
        n12328) );
  inv_1 U11813 ( .A(n12132), .Y(n12018) );
  nand2_1 U11814 ( .A(n11815), .B(n12266), .Y(n12132) );
  nand3_1 U11815 ( .A(n12208), .B(n12129), .C(n12268), .Y(n12266) );
  nand3_1 U11816 ( .A(n12270), .B(n12284), .C(n12336), .Y(n11815) );
  inv_1 U11817 ( .A(n11885), .Y(n12175) );
  nand2_1 U11818 ( .A(n12056), .B(n11941), .Y(n11885) );
  nand2_1 U11819 ( .A(n12314), .B(n12384), .Y(n11941) );
  and3_1 U11820 ( .A(n12337), .B(n12338), .C(n12287), .X(n12314) );
  nand3_1 U11821 ( .A(n12339), .B(n12341), .C(n12342), .Y(n12056) );
  nand4_1 U11822 ( .A(n11985), .B(n11956), .C(n12154), .D(n12027), .Y(n12327)
         );
  nand3_1 U11823 ( .A(n12337), .B(n12280), .C(n12343), .Y(n12027) );
  nand4_1 U11824 ( .A(n12336), .B(n12128), .C(n12084), .D(n12384), .Y(n12154)
         );
  nand4_1 U11825 ( .A(n12337), .B(n11958), .C(n11820), .D(n12384), .Y(n11956)
         );
  nand4_1 U11826 ( .A(n11822), .B(n12275), .C(n11802), .D(n12384), .Y(n11985)
         );
  nor3_1 U11827 ( .A(n12344), .B(n12030), .C(n12064), .Y(n12325) );
  nand4_1 U11828 ( .A(n12103), .B(n11793), .C(n12345), .D(n12347), .Y(n12064)
         );
  a222oi_1 U11829 ( .A1(n11986), .A2(n11900), .B1(n11858), .B2(n11870), .C1(
        n12176), .C2(n11905), .Y(n12347) );
  inv_1 U11830 ( .A(n11936), .Y(n12176) );
  nand3_1 U11831 ( .A(n12342), .B(n12348), .C(n12267), .Y(n11936) );
  inv_1 U11832 ( .A(n11935), .Y(n11858) );
  nor2_1 U11833 ( .A(n11790), .B(n11893), .Y(n11935) );
  and4_1 U11834 ( .A(n12298), .B(n12267), .C(n11820), .D(n12384), .X(n11893)
         );
  inv_1 U11835 ( .A(n12193), .Y(n11790) );
  nand3_1 U11836 ( .A(n12322), .B(n12288), .C(n11822), .Y(n12193) );
  inv_1 U11837 ( .A(n12142), .Y(n11986) );
  nand3_1 U11838 ( .A(n12276), .B(n12322), .C(n12298), .Y(n12142) );
  a21oi_1 U11839 ( .A1(n11827), .A2(n12251), .B1(n11869), .Y(n12345) );
  inv_1 U11840 ( .A(n11942), .Y(n11869) );
  nand4_1 U11841 ( .A(n11808), .B(n12296), .C(n12341), .D(n11801), .Y(n11942)
         );
  nand2_1 U11842 ( .A(n12037), .B(n12035), .Y(n12251) );
  nand3_1 U11843 ( .A(n11821), .B(n12275), .C(n12274), .Y(n12035) );
  nand3_1 U11844 ( .A(n12221), .B(n11821), .C(n11804), .Y(n12037) );
  nand2_1 U11845 ( .A(n12203), .B(n11900), .Y(n11793) );
  inv_1 U11846 ( .A(n12321), .Y(n12203) );
  nand3_1 U11847 ( .A(n12329), .B(n12275), .C(n12317), .Y(n12321) );
  nand4_1 U11848 ( .A(n12298), .B(n12287), .C(n12339), .D(n11801), .Y(n12103)
         );
  o22ai_1 U11849 ( .A1(n11838), .A2(n11901), .B1(n11884), .B2(n12281), .Y(
        n12030) );
  nand2_1 U11850 ( .A(n12268), .B(n12279), .Y(n12281) );
  and3_1 U11851 ( .A(n12349), .B(n12384), .C(n12208), .X(n12279) );
  inv_1 U11852 ( .A(n11900), .Y(n11838) );
  o21ai_0 U11853 ( .A1(n11829), .A2(n12206), .B1(n11860), .Y(n12344) );
  nor3_1 U11854 ( .A(n12145), .B(n12350), .C(n12352), .Y(n11860) );
  nand4_1 U11855 ( .A(n12106), .B(n12307), .C(n11974), .D(n12178), .Y(n12352)
         );
  or2_0 U11856 ( .A(n11794), .B(n11900), .X(n12178) );
  nand3_1 U11857 ( .A(n11803), .B(n12338), .C(n11806), .Y(n11794) );
  nand3_1 U11858 ( .A(n11808), .B(n12348), .C(n12353), .Y(n11974) );
  nor3_1 U11859 ( .A(n12356), .B(n24027), .C(n12357), .Y(n12353) );
  nand4_1 U11860 ( .A(n11988), .B(n11820), .C(n11822), .D(n11821), .Y(n12307)
         );
  nand4_1 U11861 ( .A(n11804), .B(n12311), .C(n12322), .D(n11801), .Y(n12106)
         );
  o22ai_1 U11862 ( .A1(n12190), .A2(n11805), .B1(n11953), .B2(n12048), .Y(
        n12350) );
  nand3_1 U11863 ( .A(n12358), .B(n12221), .C(n11804), .Y(n12048) );
  inv_1 U11864 ( .A(n12359), .Y(n11804) );
  nand3_1 U11865 ( .A(n11807), .B(n12317), .C(n12274), .Y(n12190) );
  nand4_1 U11866 ( .A(n12093), .B(n12309), .C(n12256), .D(n12360), .Y(n12145)
         );
  nor3_1 U11867 ( .A(n12361), .B(n12260), .C(n12051), .Y(n12360) );
  inv_1 U11868 ( .A(n12111), .Y(n12051) );
  nand4_1 U11869 ( .A(n11802), .B(n11801), .C(n11803), .D(n12362), .Y(n12111)
         );
  nor2_1 U11870 ( .A(n11819), .B(n12359), .Y(n12362) );
  and4_1 U11871 ( .A(n12294), .B(n11812), .C(n11821), .D(n12322), .X(n12260)
         );
  a21oi_1 U11872 ( .A1(n12363), .A2(n12109), .B1(n11870), .Y(n12361) );
  nand3_1 U11873 ( .A(n12238), .B(n12285), .C(n12311), .Y(n12109) );
  inv_1 U11874 ( .A(n12072), .Y(n12363) );
  o21ai_0 U11875 ( .A1(n12364), .A2(n12100), .B1(n12002), .Y(n12072) );
  nand4_1 U11876 ( .A(n12311), .B(n12238), .C(n12300), .D(n12384), .Y(n12002)
         );
  inv_1 U11877 ( .A(n12365), .Y(n12300) );
  nand3_1 U11878 ( .A(n12301), .B(n12384), .C(n11808), .Y(n12100) );
  nor2_1 U11879 ( .A(n12315), .B(n11807), .Y(n12364) );
  a22oi_1 U11880 ( .A1(n11819), .A2(n12107), .B1(n12000), .B2(n11812), .Y(
        n12256) );
  o32ai_1 U11881 ( .A1(n12366), .A2(n12367), .A3(n12365), .B1(n12368), .B2(
        n12369), .Y(n12000) );
  nand2_1 U11882 ( .A(n12267), .B(n11803), .Y(n12369) );
  nand3_1 U11883 ( .A(n12223), .B(n11801), .C(n12222), .Y(n12368) );
  inv_1 U11884 ( .A(n11806), .Y(n12367) );
  inv_1 U11885 ( .A(n12286), .Y(n12366) );
  inv_1 U11886 ( .A(n11970), .Y(n12107) );
  nand3_1 U11887 ( .A(n12296), .B(n12343), .C(n12298), .Y(n11970) );
  nor3_1 U11888 ( .A(n12370), .B(n12384), .C(n12374), .Y(n12343) );
  nand2_1 U11889 ( .A(n11818), .B(n11988), .Y(n12309) );
  inv_1 U11890 ( .A(n11819), .Y(n11988) );
  and3_1 U11891 ( .A(n12311), .B(n12286), .C(n12220), .X(n11818) );
  a21oi_1 U11892 ( .A1(n11827), .A2(n12236), .B1(n12228), .Y(n12093) );
  inv_1 U11893 ( .A(n12070), .Y(n12228) );
  nand3_1 U11894 ( .A(n12283), .B(n11821), .C(n12221), .Y(n12070) );
  and3_1 U11895 ( .A(n12329), .B(n12322), .C(n11806), .X(n12236) );
  nand2_1 U11896 ( .A(n12269), .B(n12084), .Y(n12206) );
  nor4_1 U11897 ( .A(n12252), .B(n12253), .C(n12304), .D(n12375), .Y(n12324)
         );
  mux2i_1 U11898 ( .A0(n11878), .A1(n12014), .S(n11827), .Y(n12375) );
  nand3_1 U11899 ( .A(n12323), .B(n12322), .C(n12336), .Y(n12014) );
  nand3_1 U11900 ( .A(n12329), .B(n11803), .C(n12317), .Y(n11878) );
  and2_0 U11901 ( .A(n12377), .B(n12384), .X(n12317) );
  nand4_1 U11902 ( .A(n12378), .B(n12379), .C(n12381), .D(n12382), .Y(n12304)
         );
  nor4_1 U11903 ( .A(n12259), .B(n12058), .C(n11791), .D(n12116), .Y(n12382)
         );
  inv_1 U11904 ( .A(n12141), .Y(n12116) );
  nand3_1 U11905 ( .A(n11822), .B(n11821), .C(n12286), .Y(n12141) );
  inv_1 U11906 ( .A(n11899), .Y(n11791) );
  nand4_1 U11907 ( .A(n11822), .B(n11807), .C(n11802), .D(n11801), .Y(n11899)
         );
  nor3_1 U11908 ( .A(n12383), .B(n24031), .C(n12385), .Y(n11802) );
  nor2_1 U11909 ( .A(n11830), .B(n11880), .Y(n12058) );
  nand2_1 U11910 ( .A(n12267), .B(n11957), .Y(n11830) );
  and3_1 U11911 ( .A(n12128), .B(n11801), .C(n12348), .X(n11957) );
  inv_1 U11912 ( .A(n11809), .Y(n12259) );
  nand4_1 U11913 ( .A(n12283), .B(n12377), .C(n12322), .D(n11801), .Y(n11809)
         );
  a221oi_1 U11914 ( .A1(n12248), .A2(n11819), .B1(n12250), .B2(n11953), .C1(
        n12386), .Y(n12381) );
  o22ai_1 U11915 ( .A1(n11880), .A2(n11928), .B1(n11900), .B2(n12033), .Y(
        n12386) );
  nand3_1 U11916 ( .A(n12284), .B(n12349), .C(n12270), .Y(n12033) );
  nor4_1 U11917 ( .A(n10610), .B(n12387), .C(n24024), .D(n24030), .Y(n12349)
         );
  nand2_1 U11918 ( .A(n12130), .B(n12269), .Y(n11928) );
  and2_0 U11919 ( .A(n12286), .B(n12129), .X(n12269) );
  inv_1 U11920 ( .A(n11829), .Y(n11880) );
  nand3_1 U11921 ( .A(inData[7]), .B(inData[30]), .C(inData[9]), .Y(n11829) );
  inv_1 U11922 ( .A(n12081), .Y(n12250) );
  nand3_1 U11923 ( .A(n12283), .B(n12208), .C(n12284), .Y(n12081) );
  nor2_1 U11924 ( .A(n12101), .B(n12384), .Y(n12284) );
  nand3_1 U11925 ( .A(n11134), .B(n12389), .C(inData[7]), .Y(n11819) );
  inv_1 U11926 ( .A(n11965), .Y(n12248) );
  nand3_1 U11927 ( .A(n12276), .B(n12390), .C(n12395), .Y(n11965) );
  nor3_1 U11928 ( .A(n12396), .B(n12397), .C(n12334), .Y(n12395) );
  nor3_1 U11929 ( .A(n12398), .B(n12399), .C(n11927), .Y(n12379) );
  o21ai_0 U11930 ( .A1(n11900), .A2(n12219), .B1(n11984), .Y(n11927) );
  nand2_1 U11931 ( .A(n12348), .B(n12400), .Y(n11984) );
  nor3_1 U11932 ( .A(n24025), .B(n24031), .C(n12385), .Y(n12348) );
  nand3_1 U11933 ( .A(n12285), .B(n12377), .C(n12238), .Y(n12219) );
  inv_1 U11934 ( .A(n12076), .Y(n12399) );
  a21oi_1 U11935 ( .A1(n11827), .A2(n12161), .B1(n12162), .Y(n12076) );
  and3_1 U11936 ( .A(n12311), .B(n12275), .C(n12220), .X(n12162) );
  inv_1 U11937 ( .A(n11843), .Y(n12220) );
  nand2_1 U11938 ( .A(n12329), .B(n11801), .Y(n11843) );
  nor2_1 U11939 ( .A(n12403), .B(n12404), .Y(n12311) );
  inv_1 U11940 ( .A(n11828), .Y(n12161) );
  nand3_1 U11941 ( .A(n12358), .B(n12275), .C(n12294), .Y(n11828) );
  nor3_1 U11942 ( .A(n12405), .B(n12406), .C(n12407), .Y(n12275) );
  nor3_1 U11943 ( .A(n12403), .B(n11801), .C(n12409), .Y(n12358) );
  inv_1 U11944 ( .A(n11953), .Y(n11827) );
  o21ai_0 U11945 ( .A1(n11814), .A2(n12189), .B1(n12149), .Y(n12398) );
  a22oi_1 U11946 ( .A1(n11905), .A2(n11873), .B1(n11884), .B2(n12078), .Y(
        n12149) );
  inv_1 U11947 ( .A(n11877), .Y(n12078) );
  nand3_1 U11948 ( .A(n12209), .B(n12239), .C(n12130), .Y(n11877) );
  nor3_1 U11949 ( .A(n12397), .B(n12384), .C(n12357), .Y(n12209) );
  and3_1 U11950 ( .A(n12285), .B(n12128), .C(n12130), .X(n11873) );
  nor4_1 U11951 ( .A(n12403), .B(n12410), .C(n24025), .D(n24031), .Y(n12130)
         );
  nor3_1 U11952 ( .A(n12411), .B(n24026), .C(n12407), .Y(n12128) );
  nand3_1 U11953 ( .A(n12287), .B(n11958), .C(n12323), .Y(n12189) );
  and3_1 U11954 ( .A(n12086), .B(n12257), .C(n12198), .X(n12378) );
  inv_1 U11955 ( .A(n12254), .Y(n12198) );
  o21ai_0 U11956 ( .A1(n11805), .A2(n11795), .B1(n11983), .Y(n12254) );
  nand4_1 U11957 ( .A(n11808), .B(n11884), .C(n11807), .D(n11806), .Y(n11983)
         );
  nor3_1 U11958 ( .A(n12403), .B(n12384), .C(n12409), .Y(n11806) );
  nor2_1 U11959 ( .A(n12415), .B(n12407), .Y(n11807) );
  inv_1 U11960 ( .A(n11805), .Y(n11884) );
  nor2_1 U11961 ( .A(n12374), .B(n12416), .Y(n11808) );
  nand4_1 U11962 ( .A(n12329), .B(n12301), .C(n11803), .D(n12384), .Y(n11795)
         );
  inv_1 U11963 ( .A(n12417), .Y(n12257) );
  o221ai_1 U11964 ( .A1(n11812), .A2(n12181), .B1(n11814), .B2(n12019), .C1(
        n12191), .Y(n12417) );
  nand4_1 U11965 ( .A(n12301), .B(n11801), .C(n11820), .D(n12418), .Y(n12191)
         );
  nor2_1 U11966 ( .A(n11900), .B(n12365), .Y(n12418) );
  nand2_1 U11967 ( .A(n12419), .B(n24024), .Y(n12365) );
  nand3_1 U11968 ( .A(n12342), .B(n11958), .C(n12337), .Y(n12019) );
  nor3_1 U11969 ( .A(n12356), .B(n12357), .C(n12407), .Y(n12342) );
  inv_1 U11970 ( .A(n11905), .Y(n11814) );
  nand3_1 U11971 ( .A(inData[30]), .B(n12389), .C(inData[7]), .Y(n11905) );
  nand2_1 U11972 ( .A(n12400), .B(n12341), .Y(n12181) );
  and3_1 U11973 ( .A(n12339), .B(n11801), .C(n12280), .X(n12400) );
  inv_1 U11974 ( .A(n11870), .Y(n11812) );
  nor4_1 U11975 ( .A(n11971), .B(n12080), .C(n11982), .D(n12420), .Y(n12086)
         );
  o22ai_1 U11976 ( .A1(n11900), .A2(n11898), .B1(n12192), .B2(n11953), .Y(
        n12420) );
  nand3_1 U11977 ( .A(n12303), .B(n12389), .C(n11134), .Y(n11953) );
  nand4_1 U11978 ( .A(n12221), .B(n12285), .C(n12222), .D(n12223), .Y(n12192)
         );
  and2_0 U11979 ( .A(n12283), .B(n12384), .X(n12285) );
  nor2_1 U11980 ( .A(n12415), .B(n24027), .Y(n12221) );
  nand3_1 U11981 ( .A(n11803), .B(n12338), .C(n11821), .Y(n11898) );
  nor2_1 U11982 ( .A(n12405), .B(n12397), .Y(n11803) );
  nand3_1 U11983 ( .A(inData[7]), .B(n11134), .C(inData[9]), .Y(n11900) );
  inv_1 U11984 ( .A(n11929), .Y(n11982) );
  nand3_1 U11985 ( .A(n12268), .B(n11821), .C(n12283), .Y(n11929) );
  and3_1 U11986 ( .A(n12421), .B(n11801), .C(n12422), .X(n11821) );
  nor3_1 U11987 ( .A(n24026), .B(n24027), .C(n12423), .Y(n12268) );
  inv_1 U11988 ( .A(n11990), .Y(n12080) );
  nand4_1 U11989 ( .A(n12296), .B(n12337), .C(n11822), .D(n11801), .Y(n11990)
         );
  inv_1 U11990 ( .A(n11894), .Y(n11971) );
  nand4_1 U11991 ( .A(n12287), .B(n12337), .C(n11958), .D(n11801), .Y(n11894)
         );
  nor2_1 U11992 ( .A(n12424), .B(n24025), .Y(n12337) );
  nor2_1 U11993 ( .A(n12425), .B(n12407), .Y(n12287) );
  nand2_1 U11994 ( .A(n12427), .B(n11895), .Y(n12253) );
  nand2_1 U11995 ( .A(n12125), .B(n11870), .Y(n11895) );
  nand3_1 U11996 ( .A(n11134), .B(n12303), .C(inData[9]), .Y(n11870) );
  inv_1 U11997 ( .A(n12117), .Y(n12125) );
  nand3_1 U11998 ( .A(n12084), .B(n12280), .C(n12129), .Y(n12117) );
  nor4_1 U11999 ( .A(n12383), .B(n24023), .C(n24031), .D(n24035), .Y(n12084)
         );
  mux2_1 U12000 ( .A0(n12061), .A1(n12197), .S(n11805), .X(n12427) );
  nand3_1 U12001 ( .A(n12303), .B(n12389), .C(inData[30]), .Y(n11805) );
  nand4_1 U12002 ( .A(n12286), .B(n12274), .C(n12301), .D(n11801), .Y(n12197)
         );
  nor3_1 U12003 ( .A(n10610), .B(n24024), .C(n12428), .Y(n12274) );
  nor3_1 U12004 ( .A(n12423), .B(n24026), .C(n12407), .Y(n12286) );
  nand4_1 U12005 ( .A(n12238), .B(n12208), .C(n12239), .D(n11801), .Y(n12061)
         );
  and2_0 U12006 ( .A(n12422), .B(n12223), .X(n12208) );
  and2_0 U12007 ( .A(n12431), .B(n12407), .X(n12238) );
  nand4_1 U12008 ( .A(n11910), .B(n12091), .C(n11961), .D(n12271), .Y(n12252)
         );
  nand3_1 U12009 ( .A(n12276), .B(n12341), .C(n12296), .Y(n12271) );
  nor2_1 U12010 ( .A(n12425), .B(n24027), .Y(n12296) );
  nand3_1 U12011 ( .A(n12322), .B(n12341), .C(n12276), .Y(n11961) );
  nand3_1 U12012 ( .A(n11958), .B(n11820), .C(n12323), .Y(n12091) );
  nor3_1 U12013 ( .A(n12334), .B(n11801), .C(n12396), .Y(n12323) );
  nor3_1 U12014 ( .A(n12423), .B(n12406), .C(n12407), .Y(n11820) );
  nor3_1 U12015 ( .A(n24024), .B(n24029), .C(n12428), .Y(n11958) );
  inv_1 U12016 ( .A(n11841), .Y(n11910) );
  nand2_1 U12017 ( .A(n11876), .B(n12126), .Y(n11841) );
  nand3_1 U12018 ( .A(n12129), .B(n12280), .C(n12270), .Y(n12126) );
  nor4_1 U12019 ( .A(n12403), .B(n12383), .C(n24031), .D(n24035), .Y(n12270)
         );
  nor3_1 U12020 ( .A(n24026), .B(n24027), .C(n12411), .Y(n12280) );
  and2_0 U12021 ( .A(n12239), .B(n12384), .X(n12129) );
  nor4_1 U12022 ( .A(n12387), .B(n24024), .C(n24029), .D(n24030), .Y(n12239)
         );
  nand3_1 U12023 ( .A(n12301), .B(n12276), .C(n12315), .Y(n11876) );
  inv_1 U12024 ( .A(n12101), .Y(n12315) );
  nand2_1 U12025 ( .A(n24027), .B(n12431), .Y(n12101) );
  nor3_1 U12026 ( .A(n11801), .B(n12370), .C(n12374), .Y(n12276) );
  nand2_1 U12027 ( .A(n23922), .B(n12432), .Y(n10485) );
  xnor2_1 U12028 ( .A(n12433), .B(n12434), .Y(n12432) );
  nand2_1 U12029 ( .A(n12435), .B(n12436), .Y(n12433) );
  inv_1 U12030 ( .A(n12437), .Y(n12435) );
  nand2_1 U12031 ( .A(n12438), .B(n23922), .Y(n10484) );
  xor2_1 U12032 ( .A(n12439), .B(n12443), .X(n12438) );
  xor2_1 U12033 ( .A(n12444), .B(n1144), .X(n12439) );
  o32ai_1 U12034 ( .A1(n11355), .A2(n12447), .A3(n10922), .B1(n10924), .B2(
        n12448), .Y(n10483) );
  xor2_1 U12035 ( .A(n12449), .B(n12453), .X(n12448) );
  xor2_1 U12036 ( .A(n12454), .B(n12455), .X(n12453) );
  nand4_1 U12037 ( .A(n12456), .B(n12457), .C(n12458), .D(n12459), .Y(n10482)
         );
  nand4_1 U12038 ( .A(n12460), .B(n12461), .C(n12462), .D(n10826), .Y(n12457)
         );
  or3_1 U12039 ( .A(n12463), .B(n12465), .C(n12466), .X(n12456) );
  nand2_1 U12040 ( .A(n23922), .B(n12468), .Y(n10481) );
  xor2_1 U12041 ( .A(n12469), .B(n12470), .X(n12468) );
  nor2_1 U12042 ( .A(n12471), .B(n10774), .Y(n10480) );
  xor2_1 U12043 ( .A(n12474), .B(n12477), .X(n12471) );
  xor2_1 U12044 ( .A(n12483), .B(n11525), .X(n12477) );
  xor2_1 U12045 ( .A(n12488), .B(n12489), .X(n12474) );
  nand2_1 U12046 ( .A(n12490), .B(n11500), .Y(n10479) );
  mux2_1 U12047 ( .A0(n12491), .A1(n23672), .S(n11306), .X(n12490) );
  nor2_1 U12048 ( .A(n12402), .B(n11330), .Y(n12491) );
  nand2_1 U12049 ( .A(n23922), .B(n12492), .Y(n10478) );
  xor2_1 U12050 ( .A(n12493), .B(n12494), .X(n12492) );
  xor2_1 U12051 ( .A(n12495), .B(n12496), .X(n12494) );
  xor2_1 U12052 ( .A(n12497), .B(n12297), .X(n12493) );
  o22ai_1 U12053 ( .A1(n56), .A2(n11357), .B1(n11304), .B2(n12498), .Y(n10477)
         );
  xor2_1 U12054 ( .A(outData[12]), .B(n12413), .X(n12498) );
  nor2_1 U12055 ( .A(n10774), .B(n12499), .Y(n10476) );
  xor2_1 U12056 ( .A(n12500), .B(n12501), .X(n12499) );
  nand2_1 U12057 ( .A(n12502), .B(n12503), .Y(n12501) );
  o32ai_1 U12058 ( .A1(n12504), .A2(n11150), .A3(n12505), .B1(n12507), .B2(
        n11152), .Y(n10475) );
  xor2_1 U12059 ( .A(n12508), .B(n12509), .X(n12507) );
  xor2_1 U12060 ( .A(n12512), .B(n12514), .X(n12509) );
  xor2_1 U12061 ( .A(n11197), .B(n12297), .X(n12514) );
  xor2_1 U12062 ( .A(n12519), .B(n12523), .X(n12508) );
  xor2_1 U12063 ( .A(n23932), .B(n12376), .X(n12504) );
  nor2_1 U12064 ( .A(n10774), .B(n12524), .Y(n10474) );
  xor2_1 U12065 ( .A(n12525), .B(n12526), .X(n12524) );
  xor2_1 U12066 ( .A(n12527), .B(n12528), .X(n12526) );
  xor2_1 U12067 ( .A(n12529), .B(n12530), .X(n12525) );
  nand2_1 U12068 ( .A(n12531), .B(n11500), .Y(n10473) );
  mux2_1 U12069 ( .A0(n12532), .A1(n23671), .S(n11306), .X(n12531) );
  xor2_1 U12070 ( .A(n12533), .B(n12534), .X(n12532) );
  nand2_1 U12071 ( .A(outData[10]), .B(outData[8]), .Y(n12534) );
  nor2_1 U12072 ( .A(n10774), .B(n12535), .Y(n10472) );
  xor2_1 U12073 ( .A(n12536), .B(n12537), .X(n12535) );
  xnor2_1 U12074 ( .A(n12538), .B(n12539), .Y(n12537) );
  mux2i_1 U12075 ( .A0(n61), .A1(n12540), .S(n11170), .Y(n10471) );
  nor3_1 U12076 ( .A(n11330), .B(n12346), .C(n11226), .Y(n12540) );
  o22ai_1 U12077 ( .A1(n30), .A2(n11170), .B1(n11177), .B2(n12541), .Y(n10470)
         );
  xor2_1 U12078 ( .A(n12542), .B(n12543), .X(n12541) );
  nor2_1 U12079 ( .A(n12310), .B(n11225), .Y(n12542) );
  or2_0 U12080 ( .A(n12545), .B(n12548), .X(n11170) );
  a21oi_1 U12081 ( .A1(n12550), .A2(n12551), .B1(n11304), .Y(n12545) );
  nor2_1 U12082 ( .A(n12552), .B(n11618), .Y(n11304) );
  nand2_1 U12083 ( .A(n12553), .B(n11390), .Y(n10469) );
  mux2i_1 U12084 ( .A0(n12554), .A1(n12555), .S(n11393), .Y(n12553) );
  or2_0 U12085 ( .A(n11545), .B(n756), .X(n12555) );
  o22ai_1 U12086 ( .A1(n12556), .A2(n12557), .B1(n12559), .B2(n12560), .Y(
        n12554) );
  inv_1 U12087 ( .A(n12561), .Y(n12559) );
  and2_0 U12088 ( .A(n12561), .B(n12562), .X(n12556) );
  nand4_1 U12089 ( .A(n12563), .B(n12565), .C(n12566), .D(n12567), .Y(n10468)
         );
  nand3_1 U12090 ( .A(n12568), .B(n11394), .C(n12569), .Y(n12567) );
  or3_1 U12091 ( .A(n12570), .B(n12571), .C(n12572), .X(n12566) );
  nand2_1 U12092 ( .A(n12573), .B(n12574), .Y(n12565) );
  inv_1 U12093 ( .A(n12575), .Y(n12563) );
  nand4_1 U12094 ( .A(n12576), .B(n12577), .C(n12578), .D(n12585), .Y(n10467)
         );
  nor3_1 U12095 ( .A(n12588), .B(n12589), .C(n12590), .Y(n12585) );
  a21oi_1 U12096 ( .A1(n12591), .A2(n12592), .B1(n12593), .Y(n12590) );
  a21oi_1 U12097 ( .A1(n12594), .A2(n12595), .B1(n12596), .Y(n12589) );
  a21oi_1 U12098 ( .A1(n12597), .A2(n12598), .B1(n12599), .Y(n12588) );
  nor4_1 U12099 ( .A(n12600), .B(n12601), .C(n12602), .D(n12603), .Y(n12598)
         );
  nand3_1 U12100 ( .A(n12604), .B(n12605), .C(n12606), .Y(n12600) );
  nor4_1 U12101 ( .A(n12607), .B(n12608), .C(n12609), .D(n12610), .Y(n12597)
         );
  nand3_1 U12102 ( .A(n12611), .B(n12612), .C(n12613), .Y(n12607) );
  a222oi_1 U12103 ( .A1(n12614), .A2(n12615), .B1(n12616), .B2(n12617), .C1(
        n12618), .C2(n12619), .Y(n12578) );
  inv_1 U12104 ( .A(n12620), .Y(n12614) );
  nor3_1 U12105 ( .A(n12621), .B(n12622), .C(n12623), .Y(n12577) );
  and3_1 U12106 ( .A(n12624), .B(n12625), .C(n12626), .X(n12576) );
  nor2_1 U12107 ( .A(n12627), .B(n12628), .Y(n10466) );
  xor2_1 U12108 ( .A(n12629), .B(n12630), .X(n12627) );
  xor2_1 U12109 ( .A(n12631), .B(n12632), .X(n12630) );
  nand2_1 U12110 ( .A(n12633), .B(n12634), .Y(n12631) );
  inv_1 U12111 ( .A(n12635), .Y(n12634) );
  nand2_1 U12112 ( .A(n12636), .B(n12637), .Y(n10465) );
  xor2_1 U12113 ( .A(n12638), .B(n12639), .X(n12637) );
  xor2_1 U12114 ( .A(n12640), .B(n23831), .X(n12639) );
  nand2_1 U12115 ( .A(n12641), .B(n11032), .Y(n10464) );
  mux2i_1 U12116 ( .A0(n12642), .A1(n12643), .S(n11035), .Y(n12641) );
  nand2_1 U12117 ( .A(inData[26]), .B(n12644), .Y(n12643) );
  xor2_1 U12118 ( .A(n12645), .B(n12646), .X(n12642) );
  xnor2_1 U12119 ( .A(n12647), .B(n12648), .Y(n12646) );
  xor2_1 U12120 ( .A(n12649), .B(n12650), .X(n12645) );
  nand2_1 U12121 ( .A(n12651), .B(n12652), .Y(n10463) );
  mux2i_1 U12122 ( .A0(n12653), .A1(n12654), .S(n12655), .Y(n12651) );
  xor2_1 U12123 ( .A(n12656), .B(n12657), .X(n12654) );
  nand2_1 U12124 ( .A(n18), .B(n12644), .Y(n12657) );
  inv_1 U12125 ( .A(n12430), .Y(n12644) );
  xor2_1 U12126 ( .A(n12658), .B(n12659), .X(n12653) );
  o32ai_1 U12127 ( .A1(n12660), .A2(n12661), .A3(n10678), .B1(n12662), .B2(
        n12663), .Y(n10462) );
  xor2_1 U12128 ( .A(n12664), .B(n12665), .X(n12662) );
  xor2_1 U12129 ( .A(n12666), .B(n12667), .X(n12664) );
  xor2_1 U12130 ( .A(n12668), .B(n12669), .X(n12661) );
  xor2_1 U12131 ( .A(n23856), .B(n23789), .X(n12669) );
  or2_0 U12132 ( .A(n10641), .B(n23714), .X(n12668) );
  o22ai_1 U12133 ( .A1(n10641), .A2(n12660), .B1(n12663), .B2(n12670), .Y(
        n10461) );
  xor2_1 U12134 ( .A(n12671), .B(n12672), .X(n12670) );
  xor2_1 U12135 ( .A(n12673), .B(n12430), .X(n12672) );
  o22ai_1 U12136 ( .A1(n12663), .A2(n12674), .B1(n12660), .B2(n12675), .Y(
        n10460) );
  xor2_1 U12137 ( .A(n23789), .B(n23714), .X(n12675) );
  xor2_1 U12138 ( .A(n12676), .B(n12677), .X(n12674) );
  xor2_1 U12139 ( .A(n12678), .B(n23711), .X(n12677) );
  mux2i_1 U12140 ( .A0(n12679), .A1(n12680), .S(n11097), .Y(n10459) );
  and3_1 U12141 ( .A(n23858), .B(n12681), .C(inData[14]), .X(n12680) );
  xor2_1 U12142 ( .A(n12682), .B(n12683), .X(n12679) );
  xor2_1 U12143 ( .A(n12684), .B(n12685), .X(n12683) );
  xor2_1 U12144 ( .A(n12686), .B(n12687), .X(n12682) );
  o22ai_1 U12145 ( .A1(n12688), .A2(n11097), .B1(n12689), .B2(n11094), .Y(
        n10458) );
  xor2_1 U12146 ( .A(n12690), .B(n23859), .X(n12689) );
  xnor2_1 U12147 ( .A(n12691), .B(n12692), .Y(n12688) );
  xor2_1 U12148 ( .A(n12693), .B(n12694), .X(n12692) );
  mux2i_1 U12149 ( .A0(n12695), .A1(n12696), .S(n11097), .Y(n10457) );
  nor3_1 U12150 ( .A(n12697), .B(n12698), .C(n12699), .Y(n12696) );
  xor2_1 U12151 ( .A(n23859), .B(n23814), .X(n12697) );
  xor2_1 U12152 ( .A(n12700), .B(n12701), .X(n12695) );
  nand2_1 U12153 ( .A(n12702), .B(n11377), .Y(n10456) );
  mux2i_1 U12154 ( .A0(n12703), .A1(n12704), .S(n11382), .Y(n12702) );
  xor2_1 U12155 ( .A(n12705), .B(n12706), .X(n12704) );
  xor2_1 U12156 ( .A(n12707), .B(n12708), .X(n12706) );
  xor2_1 U12157 ( .A(n12709), .B(n12710), .X(n12703) );
  xor2_1 U12158 ( .A(n23867), .B(n23767), .X(n12710) );
  nand2_1 U12159 ( .A(n23865), .B(n12711), .Y(n12709) );
  mux2i_1 U12160 ( .A0(n12712), .A1(n12713), .S(n11382), .Y(n10455) );
  xor2_1 U12161 ( .A(n12714), .B(n12715), .X(n12713) );
  xor2_1 U12162 ( .A(n23858), .B(n12716), .X(n12714) );
  nand2_1 U12163 ( .A(n12717), .B(n12711), .Y(n12712) );
  o22ai_1 U12164 ( .A1(n12718), .A2(n12719), .B1(n12720), .B2(n12721), .Y(
        n10454) );
  xor2_1 U12165 ( .A(n12722), .B(n12723), .X(n12720) );
  xor2_1 U12166 ( .A(n12724), .B(n12725), .X(n12723) );
  xor2_1 U12167 ( .A(n12726), .B(n23715), .X(n12722) );
  o22ai_1 U12168 ( .A1(n12721), .A2(n12727), .B1(n12728), .B2(n12719), .Y(
        n10453) );
  xor2_1 U12169 ( .A(n12718), .B(n23865), .X(n12728) );
  xor2_1 U12170 ( .A(n12729), .B(n12730), .X(n12727) );
  xor2_1 U12171 ( .A(n12731), .B(n11734), .X(n12730) );
  xor2_1 U12172 ( .A(n12510), .B(n12732), .X(n12729) );
  o22ai_1 U12173 ( .A1(n11333), .A2(n12733), .B1(n12734), .B2(n11331), .Y(
        n10452) );
  xor2_1 U12174 ( .A(n12735), .B(n54), .X(n12734) );
  xor2_1 U12175 ( .A(n12736), .B(n12737), .X(n12733) );
  o21ai_0 U12176 ( .A1(n12738), .A2(n12739), .B1(n12740), .Y(n12737) );
  o32ai_1 U12177 ( .A1(n11150), .A2(n12741), .A3(n10923), .B1(n12742), .B2(
        n11152), .Y(n10451) );
  xor2_1 U12178 ( .A(n12743), .B(n12744), .X(n12742) );
  xor2_1 U12179 ( .A(n12745), .B(n52), .X(n12743) );
  xor2_1 U12180 ( .A(n12746), .B(n23928), .X(n12741) );
  o221ai_1 U12181 ( .A1(n12747), .A2(n12748), .B1(n10683), .B2(n10697), .C1(
        n12749), .Y(n10450) );
  or3_1 U12182 ( .A(n10631), .B(n12750), .C(n12751), .X(n12749) );
  nor2_1 U12183 ( .A(n12752), .B(n12753), .Y(n12748) );
  o221ai_1 U12184 ( .A1(n12754), .A2(n12750), .B1(n12755), .B2(n10683), .C1(
        n12756), .Y(n10449) );
  nand2_1 U12185 ( .A(n12757), .B(n12758), .Y(n12756) );
  nand4_1 U12186 ( .A(n12759), .B(n12760), .C(n12761), .D(n12762), .Y(n12758)
         );
  nor4_1 U12187 ( .A(n10691), .B(n10722), .C(n12763), .D(n12764), .Y(n12762)
         );
  nor3_1 U12188 ( .A(n12765), .B(n10715), .C(n12766), .Y(n12761) );
  nor4_1 U12189 ( .A(n12767), .B(n12768), .C(n12769), .D(n12770), .Y(n12755)
         );
  nand3_1 U12190 ( .A(n12771), .B(n12772), .C(n12773), .Y(n12768) );
  nand4_1 U12191 ( .A(n12774), .B(n12775), .C(n12776), .D(n12777), .Y(n12767)
         );
  and2_0 U12192 ( .A(n12778), .B(n10710), .X(n12776) );
  nor4_1 U12193 ( .A(n12779), .B(n12780), .C(n12781), .D(n12782), .Y(n12754)
         );
  nand3_1 U12194 ( .A(n12783), .B(n10694), .C(n12784), .Y(n12779) );
  inv_1 U12195 ( .A(n12785), .Y(n12784) );
  nand2_1 U12196 ( .A(n23922), .B(n12786), .Y(n10448) );
  xor2_1 U12197 ( .A(n12787), .B(n12788), .X(n12786) );
  xor2_1 U12198 ( .A(n12789), .B(n12790), .X(n12788) );
  or2_0 U12199 ( .A(n50), .B(n11558), .X(n10447) );
  nand2_1 U12200 ( .A(n12791), .B(n11534), .Y(n10446) );
  or2_0 U12201 ( .A(n12792), .B(n11537), .X(n11534) );
  mux2i_1 U12202 ( .A0(n12793), .A1(n12794), .S(n11537), .Y(n12791) );
  inv_1 U12203 ( .A(n11333), .Y(n11537) );
  xor2_1 U12204 ( .A(n12795), .B(n12796), .X(n12794) );
  a21oi_1 U12205 ( .A1(n12797), .A2(n12798), .B1(n12799), .Y(n12796) );
  nand2_1 U12206 ( .A(n12800), .B(inData[30]), .Y(n12793) );
  xnor2_1 U12207 ( .A(n23706), .B(n23925), .Y(n12800) );
  mux2i_1 U12208 ( .A0(n12801), .A1(n12802), .S(n11470), .Y(n10445) );
  nor2_1 U12209 ( .A(n12803), .B(n11472), .Y(n12802) );
  xor2_1 U12210 ( .A(n11474), .B(n23936), .X(n12803) );
  nand2_1 U12211 ( .A(n23997), .B(n821), .Y(n11474) );
  xor2_1 U12212 ( .A(n12804), .B(n12805), .X(n12801) );
  xor2_1 U12213 ( .A(n10777), .B(n12806), .X(n12805) );
  xor2_1 U12214 ( .A(n12807), .B(n23971), .X(n12804) );
  nand2_1 U12215 ( .A(n12808), .B(n23922), .Y(n10444) );
  xor2_1 U12216 ( .A(n12809), .B(n12810), .X(n12808) );
  nand2_1 U12217 ( .A(n12811), .B(n12812), .Y(n12809) );
  inv_1 U12218 ( .A(n12813), .Y(n12812) );
  or2_0 U12219 ( .A(n44), .B(n11558), .X(n10443) );
  nand2_1 U12220 ( .A(n12814), .B(n23922), .Y(n10442) );
  xor2_1 U12221 ( .A(n12815), .B(n12816), .X(n12814) );
  xor2_1 U12222 ( .A(n12817), .B(n12818), .X(n12816) );
  nand2_1 U12223 ( .A(n12819), .B(n12820), .Y(n12818) );
  xor2_1 U12224 ( .A(n12821), .B(n12822), .X(n12819) );
  xor2_1 U12225 ( .A(n12823), .B(n12824), .X(n12815) );
  nand2_1 U12226 ( .A(n12825), .B(n11500), .Y(n10441) );
  mux2i_1 U12227 ( .A0(n12414), .A1(n51), .S(n11306), .Y(n12825) );
  inv_1 U12228 ( .A(n11357), .Y(n11306) );
  nand2_1 U12229 ( .A(n11418), .B(n11226), .Y(n11357) );
  o32ai_1 U12230 ( .A1(n12826), .A2(n12827), .A3(n11226), .B1(n11617), .B2(
        n12828), .Y(n10440) );
  xor2_1 U12231 ( .A(n12829), .B(n12830), .X(n12828) );
  xnor2_1 U12232 ( .A(n12831), .B(n12832), .Y(n12830) );
  xor2_1 U12233 ( .A(n12833), .B(n12834), .X(n12827) );
  xor2_1 U12234 ( .A(n23860), .B(n19), .X(n12834) );
  nand2_1 U12235 ( .A(n23712), .B(n12510), .Y(n12833) );
  nand2_1 U12236 ( .A(n12835), .B(n12836), .Y(n10439) );
  mux2i_1 U12237 ( .A0(n12837), .A1(n12838), .S(n11617), .Y(n12835) );
  xnor2_1 U12238 ( .A(n12839), .B(n12840), .Y(n12837) );
  o221ai_1 U12239 ( .A1(n12841), .A2(n12842), .B1(n12843), .B2(n12844), .C1(
        n12845), .Y(n10438) );
  o21ai_0 U12240 ( .A1(n12846), .A2(n11009), .B1(n12847), .Y(n12845) );
  nor3_1 U12241 ( .A(n12848), .B(n23709), .C(n12849), .Y(n12846) );
  a22oi_1 U12242 ( .A1(n12850), .A2(n11046), .B1(n12851), .B2(n10627), .Y(
        n12841) );
  nand2_1 U12243 ( .A(n12852), .B(n12853), .Y(n10437) );
  mux2i_1 U12244 ( .A0(n12854), .A1(n12855), .S(n12856), .Y(n12852) );
  xnor2_1 U12245 ( .A(n12857), .B(n12858), .Y(n12855) );
  xor2_1 U12246 ( .A(n12859), .B(n12860), .X(n12858) );
  nand2_1 U12247 ( .A(n12861), .B(inData[22]), .Y(n12854) );
  xor2_1 U12248 ( .A(n12862), .B(n11), .X(n12861) );
  o22ai_1 U12249 ( .A1(n12863), .A2(n12864), .B1(n12865), .B2(n12866), .Y(
        n10436) );
  xor2_1 U12250 ( .A(n12867), .B(n12868), .X(n12865) );
  xor2_1 U12251 ( .A(n9), .B(n10), .X(n12868) );
  nand2_1 U12252 ( .A(n11), .B(n12546), .Y(n12867) );
  xor2_1 U12253 ( .A(n12869), .B(n12870), .X(n12864) );
  nand2_1 U12254 ( .A(n12871), .B(n12872), .Y(n12870) );
  nand2_1 U12255 ( .A(n12873), .B(n11626), .Y(n10435) );
  mux2i_1 U12256 ( .A0(n12874), .A1(n12875), .S(n11629), .Y(n12873) );
  xor2_1 U12257 ( .A(n12876), .B(n12877), .X(n12875) );
  xor2_1 U12258 ( .A(n12878), .B(n12879), .X(n12877) );
  xor2_1 U12259 ( .A(n12880), .B(n12881), .X(n12876) );
  nand2_1 U12260 ( .A(n12882), .B(inData[28]), .Y(n12874) );
  xor2_1 U12261 ( .A(n10623), .B(n8), .X(n12882) );
  nand2_1 U12262 ( .A(n12883), .B(n11626), .Y(n10434) );
  or2_0 U12263 ( .A(n12884), .B(n11629), .X(n11626) );
  mux2i_1 U12264 ( .A0(n12885), .A1(n12886), .S(n11629), .Y(n12883) );
  inv_1 U12265 ( .A(n12887), .Y(n11629) );
  xor2_1 U12266 ( .A(n12888), .B(n12889), .X(n12886) );
  xor2_1 U12267 ( .A(n10), .B(n10936), .X(n12889) );
  xor2_1 U12268 ( .A(n12890), .B(n12891), .X(n12888) );
  nand2_1 U12269 ( .A(inData[30]), .B(n12892), .Y(n12885) );
  xnor2_1 U12270 ( .A(n1519), .B(n12893), .Y(n12892) );
  or2_0 U12271 ( .A(n12894), .B(n12515), .X(n12893) );
  o32ai_1 U12272 ( .A1(n12895), .A2(n12515), .A3(n12826), .B1(n12896), .B2(
        n12897), .Y(n10433) );
  xor2_1 U12273 ( .A(n12898), .B(n12899), .X(n12896) );
  xor2_1 U12274 ( .A(n12900), .B(n12901), .X(n12899) );
  xor2_1 U12275 ( .A(n12902), .B(n12297), .X(n12898) );
  o22ai_1 U12276 ( .A1(n12903), .A2(n12897), .B1(n12904), .B2(n12895), .Y(
        n10432) );
  xor2_1 U12277 ( .A(n1519), .B(n12894), .X(n12904) );
  xor2_1 U12278 ( .A(n12905), .B(n12906), .X(n12903) );
  xor2_1 U12279 ( .A(n12907), .B(n9), .X(n12905) );
  nand2_1 U12280 ( .A(n12908), .B(n11390), .Y(n10431) );
  nand2_1 U12281 ( .A(n12909), .B(n11393), .Y(n11390) );
  inv_1 U12282 ( .A(n11645), .Y(n12909) );
  o21ai_0 U12283 ( .A1(n11442), .A2(n11320), .B1(n11319), .Y(n11645) );
  mux2i_1 U12284 ( .A0(n12910), .A1(n12911), .S(n11393), .Y(n12908) );
  nand4_1 U12285 ( .A(n11321), .B(n11451), .C(n12912), .D(n12913), .Y(n11393)
         );
  a21oi_1 U12286 ( .A1(n11314), .A2(n11445), .B1(n12914), .Y(n12913) );
  o32ai_1 U12287 ( .A1(n12915), .A2(n24053), .A3(n10618), .B1(n11442), .B2(
        n11320), .Y(n12914) );
  nand2_1 U12288 ( .A(n12916), .B(n11314), .Y(n11321) );
  nand2_1 U12289 ( .A(n70), .B(inData[24]), .Y(n12911) );
  xor2_1 U12290 ( .A(n12917), .B(n12918), .X(n12910) );
  xor2_1 U12291 ( .A(n12919), .B(n12920), .X(n12918) );
  xor2_1 U12292 ( .A(n12921), .B(n12922), .X(n12917) );
  xor2_1 U12293 ( .A(n12923), .B(n12924), .X(n12922) );
  o32ai_1 U12294 ( .A1(n11086), .A2(n12925), .A3(n11400), .B1(n12926), .B2(
        n11402), .Y(n10430) );
  xor2_1 U12295 ( .A(n12927), .B(n12928), .X(n12926) );
  o21ai_0 U12296 ( .A1(n23921), .A2(n12929), .B1(n12930), .Y(n12927) );
  xor2_1 U12297 ( .A(n12931), .B(n12932), .X(n12925) );
  xor2_1 U12298 ( .A(n68), .B(n64), .X(n12932) );
  nand2_1 U12299 ( .A(n12580), .B(n23920), .Y(n12931) );
  nor2_1 U12300 ( .A(n10774), .B(n12933), .Y(n10429) );
  xor2_1 U12301 ( .A(n12934), .B(n12935), .X(n12933) );
  xor2_1 U12302 ( .A(n12936), .B(n12937), .X(n12935) );
  nor2_1 U12303 ( .A(n12938), .B(n12939), .Y(n12937) );
  xor2_1 U12304 ( .A(n12940), .B(n12941), .X(n12934) );
  xor2_1 U12305 ( .A(n12942), .B(n12806), .X(n12941) );
  nand2_1 U12306 ( .A(n12943), .B(n11500), .Y(n10428) );
  mux2_1 U12307 ( .A0(n12944), .A1(__________0_______18819), .S(n11418), .X(
        n12943) );
  nand2_1 U12308 ( .A(n12945), .B(n23922), .Y(n10427) );
  xor2_1 U12309 ( .A(n12946), .B(n11691), .X(n12945) );
  and2_0 U12310 ( .A(n12947), .B(n12948), .X(n11691) );
  xor2_1 U12311 ( .A(n10796), .B(n12949), .X(n12947) );
  nand2_1 U12312 ( .A(n12950), .B(n12951), .Y(n12949) );
  nand2_1 U12313 ( .A(n11693), .B(n11694), .Y(n12946) );
  nand2_1 U12314 ( .A(n12952), .B(n12953), .Y(n11694) );
  xor2_1 U12315 ( .A(n12954), .B(n11661), .X(n12952) );
  inv_1 U12316 ( .A(n11701), .Y(n12954) );
  xor2_1 U12317 ( .A(n12955), .B(n12956), .X(n11693) );
  nand2_1 U12318 ( .A(n12957), .B(n12958), .Y(n12955) );
  xor2_1 U12319 ( .A(n11661), .B(n11701), .X(n12957) );
  xor2_1 U12320 ( .A(n12959), .B(n12960), .X(n11701) );
  a21oi_1 U12321 ( .A1(n12961), .A2(n10826), .B1(n12962), .Y(n12960) );
  inv_1 U12322 ( .A(n12963), .Y(n12962) );
  o21ai_0 U12323 ( .A1(n10826), .A2(n12961), .B1(n12429), .Y(n12963) );
  xor2_1 U12324 ( .A(n12429), .B(n779), .X(n11661) );
  o32ai_1 U12325 ( .A1(n12964), .A2(n11703), .A3(n10923), .B1(n23667), .B2(
        n10924), .Y(n10426) );
  xor2_1 U12326 ( .A(outData[24]), .B(n12391), .X(n12964) );
  nor2_1 U12327 ( .A(n10774), .B(n12965), .Y(n10425) );
  xor2_1 U12328 ( .A(n12966), .B(n12967), .X(n12965) );
  xor2_1 U12329 ( .A(n12968), .B(n12969), .X(n12967) );
  nand2_1 U12330 ( .A(n12970), .B(n12971), .Y(n12969) );
  xor2_1 U12331 ( .A(n12972), .B(n12973), .X(n12970) );
  nand2_1 U12332 ( .A(n12974), .B(n11500), .Y(n10424) );
  mux2_1 U12333 ( .A0(n12975), .A1(__________0_______18818), .S(n11418), .X(
        n12974) );
  nor2_1 U12334 ( .A(n12976), .B(n11107), .Y(n12975) );
  xor2_1 U12335 ( .A(n12977), .B(n12978), .X(n12976) );
  nand2_1 U12336 ( .A(n12979), .B(n11593), .Y(n10423) );
  xor2_1 U12337 ( .A(n12980), .B(n12981), .X(n12979) );
  nand2_1 U12338 ( .A(n12982), .B(n12983), .Y(n12980) );
  xor2_1 U12339 ( .A(n12984), .B(n12985), .X(n12982) );
  mux2i_1 U12340 ( .A0(n12986), .A1(n12987), .S(n11418), .Y(n10422) );
  inv_1 U12341 ( .A(n10924), .Y(n11418) );
  xnor2_1 U12342 ( .A(n12988), .B(n12989), .Y(n12987) );
  xor2_1 U12343 ( .A(n12959), .B(n12990), .X(n12989) );
  nand2_1 U12344 ( .A(n12991), .B(n11080), .Y(n12990) );
  o21ai_0 U12345 ( .A1(n12992), .A2(n12993), .B1(n12994), .Y(n12988) );
  nor3_1 U12346 ( .A(n11175), .B(n16), .C(n10922), .Y(n12986) );
  nor2_1 U12347 ( .A(n10833), .B(n12995), .Y(n10421) );
  xor2_1 U12348 ( .A(n12996), .B(n12997), .X(n12995) );
  xor2_1 U12349 ( .A(n12998), .B(n12999), .X(n12997) );
  xor2_1 U12350 ( .A(n10796), .B(n23681), .X(n12996) );
  nand2_1 U12351 ( .A(n13000), .B(n12836), .Y(n10420) );
  mux2i_1 U12352 ( .A0(n13001), .A1(n23803), .S(n11617), .Y(n13000) );
  xor2_1 U12353 ( .A(n11737), .B(n11735), .X(n13001) );
  xnor2_1 U12354 ( .A(n11740), .B(n11738), .Y(n11735) );
  o22ai_1 U12355 ( .A1(n12998), .A2(n13002), .B1(n13003), .B2(n13004), .Y(
        n11738) );
  inv_1 U12356 ( .A(n23797), .Y(n13004) );
  nor2_1 U12357 ( .A(n13005), .B(n13006), .Y(n13003) );
  xnor2_1 U12358 ( .A(n13007), .B(n13008), .Y(n11740) );
  xor2_1 U12359 ( .A(n12579), .B(n13009), .X(n13008) );
  xor2_1 U12360 ( .A(n11725), .B(n11727), .X(n13007) );
  xnor2_1 U12361 ( .A(n13010), .B(n13011), .Y(n11725) );
  a21oi_1 U12362 ( .A1(outData[29]), .A2(n13012), .B1(n11747), .Y(n13011) );
  xnor2_1 U12363 ( .A(n12972), .B(n13013), .Y(n11747) );
  nor2_1 U12364 ( .A(outData[29]), .B(n13012), .Y(n13013) );
  xor2_1 U12365 ( .A(n13014), .B(n13015), .X(n11737) );
  a222oi_1 U12366 ( .A1(n11623), .A2(n12923), .B1(n13016), .B2(n13017), .C1(
        n13018), .C2(n13019), .Y(n13015) );
  inv_1 U12367 ( .A(n11624), .Y(n13018) );
  o21ai_0 U12368 ( .A1(n12923), .A2(n13020), .B1(n11624), .Y(n13017) );
  o21ai_0 U12369 ( .A1(n13021), .A2(n13022), .B1(n13023), .Y(n11624) );
  xor2_1 U12370 ( .A(n13016), .B(n13019), .X(n11623) );
  inv_1 U12371 ( .A(n13020), .Y(n13019) );
  o21ai_0 U12372 ( .A1(n13024), .A2(n11089), .B1(n13025), .Y(n13020) );
  xor2_1 U12373 ( .A(n12998), .B(n13026), .X(n13016) );
  xor2_1 U12374 ( .A(n23797), .B(n13005), .X(n13026) );
  inv_1 U12375 ( .A(n13002), .Y(n13005) );
  o21ai_0 U12376 ( .A1(n13027), .A2(n10612), .B1(n13012), .Y(n13002) );
  nand2_1 U12377 ( .A(n13027), .B(n10612), .Y(n13012) );
  o32ai_1 U12378 ( .A1(n11367), .A2(n818), .A3(n11133), .B1(n13028), .B2(
        n11117), .Y(n10419) );
  xor2_1 U12379 ( .A(n13029), .B(n13030), .X(n13028) );
  xor2_1 U12380 ( .A(n23803), .B(n13031), .X(n13030) );
  o221ai_1 U12381 ( .A1(n13032), .A2(n13033), .B1(n13034), .B2(n10730), .C1(
        n13035), .Y(n10418) );
  nand2_1 U12382 ( .A(n13036), .B(n13037), .Y(n13035) );
  o22ai_1 U12383 ( .A1(n13038), .A2(n13039), .B1(n13040), .B2(n13041), .Y(
        n13037) );
  nand4_1 U12384 ( .A(n13042), .B(n13043), .C(n13032), .D(n13044), .Y(n13041)
         );
  a221oi_1 U12385 ( .A1(n13045), .A2(n13046), .B1(n13047), .B2(n13048), .C1(
        n13049), .Y(n13044) );
  inv_1 U12386 ( .A(n13050), .Y(n13049) );
  nand4_1 U12387 ( .A(n13051), .B(n10736), .C(n13052), .D(n13053), .Y(n13040)
         );
  nor3_1 U12388 ( .A(n13054), .B(n13055), .C(n13056), .Y(n13053) );
  inv_1 U12389 ( .A(n10744), .Y(n13054) );
  nor4_1 U12390 ( .A(n13057), .B(n13058), .C(n13059), .D(n13060), .Y(n13034)
         );
  nand4_1 U12391 ( .A(n13061), .B(n13062), .C(n13063), .D(n13064), .Y(n13057)
         );
  nand2_1 U12392 ( .A(n13046), .B(n13065), .Y(n13062) );
  and4_1 U12393 ( .A(n13066), .B(n13067), .C(n13068), .D(n13069), .X(n13032)
         );
  nor4_1 U12394 ( .A(n13070), .B(n13071), .C(n13072), .D(n13073), .Y(n13069)
         );
  inv_1 U12395 ( .A(n13074), .Y(n13072) );
  nand3_1 U12396 ( .A(n10745), .B(n13075), .C(n13076), .Y(n13070) );
  nor3_1 U12397 ( .A(n13077), .B(n13078), .C(n13079), .Y(n13068) );
  nor2_1 U12398 ( .A(n13080), .B(n13081), .Y(n13066) );
  o21ai_0 U12399 ( .A1(n13082), .A2(n10729), .B1(n13083), .Y(n10417) );
  mux2i_1 U12400 ( .A0(n10735), .A1(n13084), .S(n13085), .Y(n13083) );
  nor4_1 U12401 ( .A(n13086), .B(n13087), .C(n13078), .D(n13088), .Y(n13085)
         );
  nand2_1 U12402 ( .A(n13089), .B(n13050), .Y(n13087) );
  nand4_1 U12403 ( .A(n13051), .B(n13090), .C(n13074), .D(n13091), .Y(n13086)
         );
  and4_1 U12404 ( .A(n11901), .B(n13092), .C(n10731), .D(n13082), .X(n13084)
         );
  nor2_1 U12405 ( .A(n13093), .B(n13094), .Y(n10731) );
  inv_1 U12406 ( .A(n13095), .Y(n13094) );
  and4_1 U12407 ( .A(n13096), .B(n13097), .C(n13098), .D(n13099), .X(n13082)
         );
  and4_1 U12408 ( .A(n13100), .B(n13101), .C(n12574), .D(n13102), .X(n13099)
         );
  nand3_1 U12409 ( .A(n13103), .B(n13104), .C(n13105), .Y(n10416) );
  a21oi_1 U12410 ( .A1(n13106), .A2(n11901), .B1(n13107), .Y(n13105) );
  a21oi_1 U12411 ( .A1(n13108), .A2(n13109), .B1(n13033), .Y(n13107) );
  nor4_1 U12412 ( .A(n13110), .B(n13111), .C(n13112), .D(n13113), .Y(n13109)
         );
  nand4_1 U12413 ( .A(n13075), .B(n13114), .C(n13115), .D(n13116), .Y(n13110)
         );
  nor4_1 U12414 ( .A(n13117), .B(n13118), .C(n13058), .D(n13119), .Y(n13108)
         );
  inv_1 U12415 ( .A(n13120), .Y(n13058) );
  nand3_1 U12416 ( .A(n13052), .B(n13121), .C(n13122), .Y(n13117) );
  nand4_1 U12417 ( .A(n13123), .B(n13124), .C(n13125), .D(n13126), .Y(n13106)
         );
  a211oi_1 U12418 ( .A1(n13046), .A2(n13065), .B1(n13127), .C1(n13081), .Y(
        n13126) );
  inv_1 U12419 ( .A(n13128), .Y(n13123) );
  o21ai_0 U12420 ( .A1(n13129), .A2(n13130), .B1(n13036), .Y(n13104) );
  nand4_1 U12421 ( .A(n13131), .B(n13132), .C(n13133), .D(n13134), .Y(n13130)
         );
  and3_1 U12422 ( .A(n13135), .B(n13097), .C(n13136), .X(n13134) );
  inv_1 U12423 ( .A(n13060), .Y(n13132) );
  nand4_1 U12424 ( .A(n13137), .B(n13138), .C(n13139), .D(n13140), .Y(n13060)
         );
  inv_1 U12425 ( .A(n13141), .Y(n13131) );
  nand4_1 U12426 ( .A(n10743), .B(n13142), .C(n13050), .D(n13143), .Y(n13129)
         );
  nor3_1 U12427 ( .A(n13144), .B(n13145), .C(n13146), .Y(n13143) );
  inv_1 U12428 ( .A(n13147), .Y(n13103) );
  o221ai_1 U12429 ( .A1(n10730), .A2(n13148), .B1(n13149), .B2(n13033), .C1(
        n13150), .Y(n10415) );
  a21oi_1 U12430 ( .A1(n13036), .A2(n13151), .B1(n13152), .Y(n13150) );
  nand4_1 U12431 ( .A(n13133), .B(n13042), .C(n13153), .D(n13154), .Y(n13151)
         );
  nor4_1 U12432 ( .A(n13081), .B(n13155), .C(n13156), .D(n13157), .Y(n13154)
         );
  nor2_1 U12433 ( .A(n13158), .B(n13159), .Y(n13155) );
  nor4_1 U12434 ( .A(n13160), .B(n13161), .C(n13162), .D(n13163), .Y(n13133)
         );
  o21ai_0 U12435 ( .A1(n13164), .A2(n13158), .B1(n13096), .Y(n13163) );
  nor3_1 U12436 ( .A(n13165), .B(n13166), .C(n13167), .Y(n13149) );
  inv_1 U12437 ( .A(n13168), .Y(n13166) );
  nand3_1 U12438 ( .A(n13102), .B(n13091), .C(n13097), .Y(n13165) );
  nor3_1 U12439 ( .A(n13169), .B(n13145), .C(n12599), .Y(n13148) );
  o221ai_1 U12440 ( .A1(n10730), .A2(n13170), .B1(n13171), .B2(n10729), .C1(
        n13172), .Y(n10414) );
  a21oi_1 U12441 ( .A1(n10735), .A2(n13173), .B1(n13147), .Y(n13172) );
  nand3_1 U12442 ( .A(n13174), .B(n13175), .C(n13176), .Y(n13147) );
  o21ai_0 U12443 ( .A1(n13177), .A2(n13178), .B1(n11901), .Y(n13176) );
  nand3_1 U12444 ( .A(n10735), .B(n13179), .C(n13180), .Y(n13175) );
  o21ai_0 U12445 ( .A1(n13181), .A2(n13182), .B1(n13036), .Y(n13174) );
  nand4_1 U12446 ( .A(n13183), .B(n13184), .C(n13185), .D(n13186), .Y(n13173)
         );
  nor4_1 U12447 ( .A(n13160), .B(n13187), .C(n13157), .D(n13059), .Y(n13186)
         );
  nand3_1 U12448 ( .A(n12574), .B(n13188), .C(n13189), .Y(n13059) );
  inv_1 U12449 ( .A(n10745), .Y(n13160) );
  inv_1 U12450 ( .A(n13088), .Y(n13184) );
  nand4_1 U12451 ( .A(n13190), .B(n13052), .C(n13076), .D(n13191), .Y(n13088)
         );
  nand2_1 U12452 ( .A(n13180), .B(n13048), .Y(n13190) );
  inv_1 U12453 ( .A(n13118), .Y(n13183) );
  nand3_1 U12454 ( .A(n13100), .B(n13192), .C(n13193), .Y(n13118) );
  nor4_1 U12455 ( .A(n13194), .B(n13195), .C(n13119), .D(n13196), .Y(n13171)
         );
  nand3_1 U12456 ( .A(n13197), .B(n13198), .C(n13102), .Y(n13119) );
  nand3_1 U12457 ( .A(n13199), .B(n13200), .C(n13042), .Y(n13195) );
  a22oi_1 U12458 ( .A1(n13201), .A2(n13046), .B1(n13179), .B2(n13202), .Y(
        n13042) );
  nand4_1 U12459 ( .A(n13101), .B(n13115), .C(n13139), .D(n13203), .Y(n13194)
         );
  a211oi_1 U12460 ( .A1(n13045), .A2(n13180), .B1(n13204), .C1(n13205), .Y(
        n13203) );
  a21oi_1 U12461 ( .A1(n13206), .A2(n13207), .B1(n13039), .Y(n13205) );
  nor4_1 U12462 ( .A(n13208), .B(n13209), .C(n13210), .D(n13211), .Y(n13170)
         );
  nand3_1 U12463 ( .A(n13212), .B(n13116), .C(n13213), .Y(n13209) );
  nand4_1 U12464 ( .A(n13153), .B(n13214), .C(n13215), .D(n13216), .Y(n13208)
         );
  a21oi_1 U12465 ( .A1(n13217), .A2(n13218), .B1(n10733), .Y(n13215) );
  and3_1 U12466 ( .A(n13219), .B(n13140), .C(n13220), .X(n13153) );
  o221ai_1 U12467 ( .A1(n10730), .A2(n13221), .B1(n13222), .B2(n13033), .C1(
        n13223), .Y(n10413) );
  o21ai_0 U12468 ( .A1(n13224), .A2(n13225), .B1(n13036), .Y(n13223) );
  o221ai_1 U12469 ( .A1(n13226), .A2(n13206), .B1(n13158), .B2(n13227), .C1(
        n13228), .Y(n13225) );
  or4_1 U12470 ( .A(n13146), .B(n13229), .C(n13161), .D(n13073), .X(n13224) );
  inv_1 U12471 ( .A(n13115), .Y(n13073) );
  nor3_1 U12472 ( .A(n13230), .B(n13079), .C(n13231), .Y(n13222) );
  nor4_1 U12473 ( .A(n13232), .B(n13233), .C(n13113), .D(n13127), .Y(n13221)
         );
  nand3_1 U12474 ( .A(n13234), .B(n13235), .C(n13236), .Y(n13232) );
  o21ai_0 U12475 ( .A1(n13237), .A2(n13033), .B1(n13238), .Y(n10412) );
  mux2i_1 U12476 ( .A0(n13036), .A1(n13239), .S(n13240), .Y(n13238) );
  nor4_1 U12477 ( .A(n13241), .B(n13242), .C(n13187), .D(n13243), .Y(n13240)
         );
  inv_1 U12478 ( .A(n13189), .Y(n13243) );
  nand3_1 U12479 ( .A(n13235), .B(n13213), .C(n10736), .Y(n13242) );
  nand4_1 U12480 ( .A(n13125), .B(n13098), .C(n13216), .D(n13220), .Y(n13241)
         );
  and4_1 U12481 ( .A(n13244), .B(n13245), .C(n13135), .D(n13246), .X(n13098)
         );
  nor3_1 U12482 ( .A(n13247), .B(n13161), .C(n13248), .Y(n13246) );
  nor4_1 U12483 ( .A(n13249), .B(n13250), .C(n13251), .D(n13252), .Y(n13239)
         );
  nand3_1 U12484 ( .A(n11901), .B(n13101), .C(n13219), .Y(n13250) );
  nand4_1 U12485 ( .A(n13237), .B(n13253), .C(n13193), .D(n13043), .Y(n13249)
         );
  and3_1 U12486 ( .A(n13092), .B(n13254), .C(n13255), .X(n13043) );
  a21oi_1 U12487 ( .A1(n13217), .A2(n13256), .B1(n13257), .Y(n13255) );
  inv_1 U12488 ( .A(n13199), .Y(n13257) );
  a21oi_1 U12489 ( .A1(n13258), .A2(n13259), .B1(n13144), .Y(n13199) );
  nand2_1 U12490 ( .A(n13260), .B(n13261), .Y(n13092) );
  nor4_1 U12491 ( .A(n13262), .B(n10740), .C(n13080), .D(n10733), .Y(n13261)
         );
  nand3_1 U12492 ( .A(n13263), .B(n13264), .C(n13265), .Y(n10733) );
  nand3_1 U12493 ( .A(n10736), .B(n13101), .C(n13220), .Y(n13262) );
  nor4_1 U12494 ( .A(n13266), .B(n13169), .C(n13231), .D(n13233), .Y(n13260)
         );
  nand4_1 U12495 ( .A(n13267), .B(n13268), .C(n13269), .D(n13270), .Y(n13233)
         );
  nor4_1 U12496 ( .A(n13271), .B(n13272), .C(n13111), .D(n13273), .Y(n13270)
         );
  inv_1 U12497 ( .A(n13076), .Y(n13273) );
  nand2_1 U12498 ( .A(n13274), .B(n13212), .Y(n13272) );
  inv_1 U12499 ( .A(n13090), .Y(n13271) );
  nor3_1 U12500 ( .A(n10742), .B(n13162), .C(n13177), .Y(n13269) );
  inv_1 U12501 ( .A(n13245), .Y(n13177) );
  nand3_1 U12502 ( .A(n13063), .B(n13188), .C(n13197), .Y(n10742) );
  inv_1 U12503 ( .A(n13156), .Y(n13268) );
  nand2_1 U12504 ( .A(n13100), .B(n13050), .Y(n13156) );
  nand2_1 U12505 ( .A(n13275), .B(n13276), .Y(n13050) );
  inv_1 U12506 ( .A(n13167), .Y(n13267) );
  nand4_1 U12507 ( .A(n13124), .B(n13277), .C(n13214), .D(n13278), .Y(n13167)
         );
  and4_1 U12508 ( .A(n13116), .B(n13139), .C(n10744), .D(n10743), .X(n13278)
         );
  and3_1 U12509 ( .A(n13279), .B(n13189), .C(n13280), .X(n13124) );
  nand4_1 U12510 ( .A(n13097), .B(n10745), .C(n13281), .D(n13140), .Y(n13231)
         );
  nand2_1 U12511 ( .A(n13282), .B(n13275), .Y(n10745) );
  nand4_1 U12512 ( .A(n13115), .B(n13192), .C(n13052), .D(n13283), .Y(n13169)
         );
  nor2_1 U12513 ( .A(n13093), .B(n13077), .Y(n13283) );
  nand3_1 U12514 ( .A(n13095), .B(n13234), .C(n13284), .Y(n13077) );
  nand4_1 U12515 ( .A(n13254), .B(n13064), .C(n13285), .D(n13286), .Y(n13093)
         );
  and4_1 U12516 ( .A(n13287), .B(n13288), .C(n13122), .D(n13136), .X(n13286)
         );
  nor3_1 U12517 ( .A(n13056), .B(n13289), .C(n13144), .Y(n13285) );
  inv_1 U12518 ( .A(n13290), .Y(n13144) );
  inv_1 U12519 ( .A(n13114), .Y(n13056) );
  nand3_1 U12520 ( .A(n13228), .B(n13135), .C(n13138), .Y(n13266) );
  and4_1 U12521 ( .A(n13291), .B(n13292), .C(n13293), .D(n13294), .X(n13228)
         );
  and4_1 U12522 ( .A(n13102), .B(n13200), .C(n13168), .D(n13244), .X(n13294)
         );
  nor3_1 U12523 ( .A(n13247), .B(n13081), .C(n13251), .Y(n13200) );
  inv_1 U12524 ( .A(n13295), .Y(n13081) );
  nor2_1 U12525 ( .A(n13296), .B(n13158), .Y(n13247) );
  nand2_1 U12526 ( .A(n13275), .B(n13297), .Y(n13102) );
  nor3_1 U12527 ( .A(n13298), .B(n13055), .C(n12599), .Y(n13293) );
  and4_1 U12528 ( .A(n13185), .B(n13061), .C(n13299), .D(n13300), .X(n13237)
         );
  nor4_1 U12529 ( .A(n13301), .B(n13302), .C(n13145), .D(n13303), .Y(n13300)
         );
  inv_1 U12530 ( .A(n13281), .Y(n13302) );
  nand3_1 U12531 ( .A(n13090), .B(n13277), .C(n13291), .Y(n13301) );
  and3_1 U12532 ( .A(n13067), .B(n13265), .C(n13089), .X(n13299) );
  nor4_1 U12533 ( .A(n10740), .B(n13304), .C(n13210), .D(n13182), .Y(n13067)
         );
  inv_1 U12534 ( .A(n13197), .Y(n13304) );
  nand3_1 U12535 ( .A(n13142), .B(n13198), .C(n13236), .Y(n10740) );
  and4_1 U12536 ( .A(n13075), .B(n13305), .C(n10744), .D(n13306), .X(n13185)
         );
  and2_0 U12537 ( .A(n10743), .B(n13063), .X(n13306) );
  nand3_1 U12538 ( .A(n13307), .B(n13308), .C(n13309), .Y(n10743) );
  o211ai_1 U12539 ( .A1(n13310), .A2(n13033), .B1(n13311), .C1(n13312), .Y(
        n10411) );
  a21oi_1 U12540 ( .A1(n13036), .A2(n13313), .B1(n13152), .Y(n13312) );
  o22ai_1 U12541 ( .A1(n13314), .A2(n10729), .B1(n13315), .B2(n13033), .Y(
        n13152) );
  nor2_1 U12542 ( .A(n13316), .B(n13178), .Y(n13315) );
  a211oi_1 U12543 ( .A1(n13317), .A2(n13179), .B1(n13318), .C1(n13181), .Y(
        n13314) );
  inv_1 U12544 ( .A(n10736), .Y(n13181) );
  nand2_1 U12545 ( .A(n13319), .B(n13179), .Y(n10736) );
  inv_1 U12546 ( .A(n13265), .Y(n13318) );
  nor2_1 U12547 ( .A(n13127), .B(n13146), .Y(n13265) );
  and2_0 U12548 ( .A(n13320), .B(n13297), .X(n13146) );
  and2_0 U12549 ( .A(n13276), .B(n13308), .X(n13127) );
  nand4_1 U12550 ( .A(n13321), .B(n13288), .C(n13322), .D(n13323), .Y(n13313)
         );
  nor4_1 U12551 ( .A(n13324), .B(n13141), .C(n13325), .D(n13128), .Y(n13323)
         );
  inv_1 U12552 ( .A(n13135), .Y(n13325) );
  nor3_1 U12553 ( .A(n13229), .B(n13326), .C(n13327), .Y(n13135) );
  o22ai_1 U12554 ( .A1(n13206), .A2(n13164), .B1(n13159), .B2(n13207), .Y(
        n13327) );
  a21oi_1 U12555 ( .A1(n13328), .A2(n13329), .B1(n13226), .Y(n13326) );
  a21oi_1 U12556 ( .A1(n13038), .A2(n13328), .B1(n13164), .Y(n13229) );
  nand3_1 U12557 ( .A(n10744), .B(n13101), .C(n13220), .Y(n13141) );
  o21ai_0 U12558 ( .A1(n13048), .A2(n13330), .B1(n13319), .Y(n13101) );
  nand3_1 U12559 ( .A(n13168), .B(n13122), .C(n13214), .Y(n13324) );
  inv_1 U12560 ( .A(n13252), .Y(n13214) );
  a21oi_1 U12561 ( .A1(n13202), .A2(n13045), .B1(n13331), .Y(n13168) );
  nor4_1 U12562 ( .A(n13161), .B(n13332), .C(n13298), .D(n13187), .Y(n13322)
         );
  inv_1 U12563 ( .A(n13219), .Y(n13298) );
  inv_1 U12564 ( .A(n13139), .Y(n13332) );
  nand2_1 U12565 ( .A(n13201), .B(n13180), .Y(n13139) );
  a21oi_1 U12566 ( .A1(n13038), .A2(n13207), .B1(n13039), .Y(n13161) );
  and4_1 U12567 ( .A(n13333), .B(n13334), .C(n13335), .D(n13075), .X(n13288)
         );
  nand3_1 U12568 ( .A(n13336), .B(n24013), .C(n13218), .Y(n13333) );
  a21oi_1 U12569 ( .A1(n13337), .A2(n13330), .B1(n13162), .Y(n13321) );
  inv_1 U12570 ( .A(n13051), .Y(n13162) );
  inv_1 U12571 ( .A(n10729), .Y(n13036) );
  o21ai_0 U12572 ( .A1(n13338), .A2(n13339), .B1(n11901), .Y(n13311) );
  nand4_1 U12573 ( .A(n13340), .B(n13136), .C(n13097), .D(n13295), .Y(n13339)
         );
  nand2_1 U12574 ( .A(n13317), .B(n13048), .Y(n13295) );
  inv_1 U12575 ( .A(n13159), .Y(n13048) );
  nand2_1 U12576 ( .A(n13282), .B(n13341), .Y(n13097) );
  nand4_1 U12577 ( .A(n13189), .B(n13274), .C(n13197), .D(n13236), .Y(n13338)
         );
  nand3_1 U12578 ( .A(n13307), .B(n13342), .C(n13320), .Y(n13197) );
  nand2_1 U12579 ( .A(n13046), .B(n13179), .Y(n13189) );
  nor4_1 U12580 ( .A(n13343), .B(n13344), .C(n13345), .D(n13346), .Y(n13310)
         );
  inv_1 U12581 ( .A(n13287), .Y(n13346) );
  inv_1 U12582 ( .A(n13064), .Y(n13345) );
  nand3_1 U12583 ( .A(n13115), .B(n13100), .C(n13290), .Y(n13344) );
  nand2_1 U12584 ( .A(n13180), .B(n13347), .Y(n13115) );
  nand3_1 U12585 ( .A(n13348), .B(n13216), .C(n13349), .Y(n13343) );
  and3_1 U12586 ( .A(n10738), .B(n13263), .C(n13090), .X(n13349) );
  nor2_1 U12587 ( .A(n12599), .B(n13204), .Y(n10738) );
  inv_1 U12588 ( .A(n13078), .Y(n13216) );
  nand2_1 U12589 ( .A(n13121), .B(n13279), .Y(n13078) );
  nand3_1 U12590 ( .A(n13350), .B(n13351), .C(n13309), .Y(n13279) );
  nand3_1 U12591 ( .A(n13350), .B(n13342), .C(n13307), .Y(n13121) );
  inv_1 U12592 ( .A(n13230), .Y(n13348) );
  nand4_1 U12593 ( .A(n13198), .B(n13192), .C(n13142), .D(n13352), .Y(n13230)
         );
  nor2_1 U12594 ( .A(n13080), .B(n13353), .Y(n13352) );
  inv_1 U12595 ( .A(n13052), .Y(n13353) );
  nand3_1 U12596 ( .A(n13307), .B(n13354), .C(n13320), .Y(n13052) );
  nand3_1 U12597 ( .A(n13307), .B(n13342), .C(n13341), .Y(n13198) );
  o221ai_1 U12598 ( .A1(n13355), .A2(n10730), .B1(n13356), .B2(n10729), .C1(
        n13357), .Y(n10410) );
  o21ai_0 U12599 ( .A1(n13358), .A2(n13359), .B1(n10735), .Y(n13357) );
  inv_1 U12600 ( .A(n13033), .Y(n10735) );
  nand2_1 U12601 ( .A(inData[13]), .B(n11901), .Y(n13033) );
  nand4_1 U12602 ( .A(n13193), .B(n13137), .C(n13340), .D(n13360), .Y(n13359)
         );
  nor3_1 U12603 ( .A(n13252), .B(n10741), .C(n13079), .Y(n13360) );
  o211ai_1 U12604 ( .A1(n13159), .A2(n13038), .B1(n13220), .C1(n13089), .Y(
        n13079) );
  a21oi_1 U12605 ( .A1(n13179), .A2(n13180), .B1(n13316), .Y(n13089) );
  nor2_1 U12606 ( .A(n13207), .B(n13226), .Y(n13316) );
  inv_1 U12607 ( .A(n13047), .Y(n13207) );
  nand2_1 U12608 ( .A(n13065), .B(n13202), .Y(n13220) );
  inv_1 U12609 ( .A(n13284), .Y(n10741) );
  nand2_1 U12610 ( .A(n13297), .B(n13308), .Y(n13284) );
  o21ai_0 U12611 ( .A1(n13039), .A2(n13328), .B1(n13074), .Y(n13252) );
  nand3_1 U12612 ( .A(n13354), .B(n13350), .C(n13307), .Y(n13074) );
  and3_1 U12613 ( .A(n13253), .B(n13245), .C(n13361), .X(n13340) );
  nor3_1 U12614 ( .A(n13303), .B(n13145), .C(n13289), .Y(n13361) );
  inv_1 U12615 ( .A(n13213), .Y(n13289) );
  nand2_1 U12616 ( .A(n13362), .B(n13363), .Y(n13213) );
  inv_1 U12617 ( .A(n13212), .Y(n13145) );
  nand2_1 U12618 ( .A(n13047), .B(n13179), .Y(n13212) );
  inv_1 U12619 ( .A(n13140), .Y(n13303) );
  nand2_1 U12620 ( .A(n13330), .B(n13317), .Y(n13140) );
  nand2_1 U12621 ( .A(n13297), .B(n13350), .Y(n13245) );
  and4_1 U12622 ( .A(n13076), .B(n13188), .C(n13114), .D(n13095), .X(n13253)
         );
  nand2_1 U12623 ( .A(n13364), .B(n13363), .Y(n13095) );
  nand2_1 U12624 ( .A(n13218), .B(n13258), .Y(n13114) );
  nand2_1 U12625 ( .A(n13341), .B(n13365), .Y(n13188) );
  nand3_1 U12626 ( .A(n13275), .B(n13307), .C(n13309), .Y(n13076) );
  and4_1 U12627 ( .A(n13090), .B(n13191), .C(n13219), .D(n13366), .X(n13137)
         );
  a21oi_1 U12628 ( .A1(n13045), .A2(n13202), .B1(n13187), .Y(n13366) );
  inv_1 U12629 ( .A(n13292), .Y(n13187) );
  nand2_1 U12630 ( .A(n13065), .B(n13319), .Y(n13292) );
  nand2_1 U12631 ( .A(n13065), .B(n13317), .Y(n13219) );
  nand2_1 U12632 ( .A(n13276), .B(n13320), .Y(n13191) );
  nor3_1 U12633 ( .A(n13367), .B(n13368), .C(n13369), .Y(n13276) );
  nand2_1 U12634 ( .A(n13370), .B(n13320), .Y(n13090) );
  a21oi_1 U12635 ( .A1(n13364), .A2(n13218), .B1(n13371), .Y(n13193) );
  inv_1 U12636 ( .A(n13334), .Y(n13371) );
  nand2_1 U12637 ( .A(n13258), .B(n13363), .Y(n13334) );
  nand4_1 U12638 ( .A(n13142), .B(n13075), .C(n13236), .D(n13372), .Y(n13358)
         );
  nor3_1 U12639 ( .A(n13182), .B(n13373), .C(n13055), .Y(n13372) );
  nor2_1 U12640 ( .A(n13329), .B(n13159), .Y(n13055) );
  inv_1 U12641 ( .A(n13202), .Y(n13329) );
  inv_1 U12642 ( .A(n13116), .Y(n13373) );
  nand2_1 U12643 ( .A(n13330), .B(n13047), .Y(n13116) );
  inv_1 U12644 ( .A(n13091), .Y(n13182) );
  nand3_1 U12645 ( .A(n13308), .B(n13351), .C(n13309), .Y(n13091) );
  nand2_1 U12646 ( .A(n13370), .B(n13350), .Y(n13236) );
  nand2_1 U12647 ( .A(n13259), .B(n13364), .Y(n13075) );
  nand3_1 U12648 ( .A(n13308), .B(n13354), .C(n13307), .Y(n13142) );
  nand2_1 U12649 ( .A(n13374), .B(n11901), .Y(n10729) );
  nor4_1 U12650 ( .A(n13375), .B(n13376), .C(n13112), .D(n13204), .Y(n13356)
         );
  inv_1 U12651 ( .A(n13277), .Y(n13204) );
  nand2_1 U12652 ( .A(n13370), .B(n13275), .Y(n13277) );
  inv_1 U12653 ( .A(n13264), .Y(n13112) );
  nand2_1 U12654 ( .A(n13350), .B(n13365), .Y(n13264) );
  nand3_1 U12655 ( .A(n13290), .B(n13192), .C(n10744), .Y(n13376) );
  nand2_1 U12656 ( .A(n13341), .B(n13370), .Y(n10744) );
  nor3_1 U12657 ( .A(n13368), .B(n24002), .C(n13377), .Y(n13370) );
  nand2_1 U12658 ( .A(n13045), .B(n13047), .Y(n13192) );
  nor3_1 U12659 ( .A(n13378), .B(n13379), .C(n13380), .Y(n13047) );
  inv_1 U12660 ( .A(n13164), .Y(n13045) );
  nand2_1 U12661 ( .A(n13256), .B(n13364), .Y(n13290) );
  nor2_1 U12662 ( .A(n13381), .B(n13382), .Y(n13364) );
  nand4_1 U12663 ( .A(n13244), .B(n13096), .C(n13291), .D(n13051), .Y(n13375)
         );
  nand2_1 U12664 ( .A(n13308), .B(n13365), .Y(n13051) );
  and2_0 U12665 ( .A(n13351), .B(n13342), .X(n13365) );
  and3_1 U12666 ( .A(n13383), .B(n13384), .C(n13385), .X(n13342) );
  inv_1 U12667 ( .A(n13178), .Y(n13291) );
  nor2_1 U12668 ( .A(n13206), .B(n13159), .Y(n13178) );
  nand2_1 U12669 ( .A(n13386), .B(n13387), .Y(n13159) );
  inv_1 U12670 ( .A(n13251), .Y(n13096) );
  o22ai_1 U12671 ( .A1(n13158), .A2(n13226), .B1(n13296), .B2(n13328), .Y(
        n13251) );
  inv_1 U12672 ( .A(n13388), .Y(n13244) );
  o221ai_1 U12673 ( .A1(n13389), .A2(n13206), .B1(n13158), .B2(n13164), .C1(
        n13390), .Y(n13388) );
  o21ai_0 U12674 ( .A1(n13202), .A2(n13317), .B1(n13179), .Y(n13390) );
  inv_1 U12675 ( .A(n13391), .Y(n13179) );
  inv_1 U12676 ( .A(n13319), .Y(n13158) );
  nor3_1 U12677 ( .A(n13392), .B(n13382), .C(n13380), .Y(n13319) );
  nor2_1 U12678 ( .A(n13330), .B(n13065), .Y(n13389) );
  inv_1 U12679 ( .A(n13039), .Y(n13065) );
  nand2_1 U12680 ( .A(n13386), .B(n13385), .Y(n13039) );
  inv_1 U12681 ( .A(n11901), .Y(n10730) );
  nand3_1 U12682 ( .A(n12322), .B(n12288), .C(n12339), .Y(n11901) );
  and2_0 U12683 ( .A(n12384), .B(n12341), .X(n12288) );
  nor2_1 U12684 ( .A(n12404), .B(n24023), .Y(n12341) );
  nor2_1 U12685 ( .A(n12423), .B(n12397), .Y(n12322) );
  nand2_1 U12686 ( .A(n24026), .B(n12407), .Y(n12397) );
  nor4_1 U12687 ( .A(n13393), .B(n13394), .C(n13128), .D(n13196), .Y(n13355)
         );
  nand4_1 U12688 ( .A(n13125), .B(n13061), .C(n13281), .D(n13234), .Y(n13196)
         );
  nand2_1 U12689 ( .A(n13317), .B(n13347), .Y(n13234) );
  inv_1 U12690 ( .A(n13296), .Y(n13347) );
  nand2_1 U12691 ( .A(n13330), .B(n13202), .Y(n13281) );
  nor2_1 U12692 ( .A(n13395), .B(n13380), .Y(n13202) );
  nor2_1 U12693 ( .A(n13111), .B(n13331), .Y(n13061) );
  nor2_1 U12694 ( .A(n13206), .B(n13296), .Y(n13331) );
  nand2_1 U12695 ( .A(n13396), .B(n13397), .Y(n13296) );
  nor2_1 U12696 ( .A(n13328), .B(n13227), .Y(n13111) );
  inv_1 U12697 ( .A(n13046), .Y(n13328) );
  nor3_1 U12698 ( .A(n13380), .B(n13398), .C(n13399), .Y(n13046) );
  and3_1 U12699 ( .A(n13335), .B(n13064), .C(n13287), .X(n13125) );
  nand2_1 U12700 ( .A(n13217), .B(n13363), .Y(n13287) );
  and3_1 U12701 ( .A(n13400), .B(n13397), .C(n11751), .X(n13363) );
  nand2_1 U12702 ( .A(n13217), .B(n13259), .Y(n13064) );
  nand2_1 U12703 ( .A(n13258), .B(n13256), .Y(n13335) );
  nand2_1 U12704 ( .A(n13254), .B(n13063), .Y(n13128) );
  nand2_1 U12705 ( .A(n13282), .B(n13350), .Y(n13063) );
  nor3_1 U12706 ( .A(n13401), .B(n24002), .C(n13377), .Y(n13282) );
  nand2_1 U12707 ( .A(n13218), .B(n13362), .Y(n13254) );
  nand3_1 U12708 ( .A(n13138), .B(n13136), .C(n13120), .Y(n13394) );
  a21oi_1 U12709 ( .A1(n13218), .A2(n13217), .B1(n13248), .Y(n13120) );
  inv_1 U12710 ( .A(n13274), .Y(n13248) );
  nand3_1 U12711 ( .A(n13320), .B(n13351), .C(n13309), .Y(n13274) );
  inv_1 U12712 ( .A(n13402), .Y(n13309) );
  nor2_1 U12713 ( .A(n13403), .B(n13404), .Y(n13320) );
  and2_0 U12714 ( .A(n13396), .B(n13405), .X(n13218) );
  a21oi_1 U12715 ( .A1(n13258), .A2(n13259), .B1(n13210), .Y(n13136) );
  and2_0 U12716 ( .A(n13256), .B(n13362), .X(n13210) );
  nor2_1 U12717 ( .A(n13381), .B(n13404), .Y(n13258) );
  inv_1 U12718 ( .A(n13157), .Y(n13138) );
  o21ai_0 U12719 ( .A1(n13226), .A2(n13206), .B1(n13235), .Y(n13157) );
  nand2_1 U12720 ( .A(n13201), .B(n13317), .Y(n13235) );
  nor3_1 U12721 ( .A(n13403), .B(n13382), .C(n13380), .Y(n13317) );
  inv_1 U12722 ( .A(n13226), .Y(n13201) );
  nand2_1 U12723 ( .A(n13396), .B(n13386), .Y(n13226) );
  nand3_1 U12724 ( .A(n13122), .B(n13280), .C(n13406), .Y(n13393) );
  nor3_1 U12725 ( .A(n13080), .B(n13407), .C(n13113), .Y(n13406) );
  inv_1 U12726 ( .A(n13263), .Y(n13113) );
  nand3_1 U12727 ( .A(n13354), .B(n13351), .C(n13308), .Y(n13263) );
  inv_1 U12728 ( .A(n13100), .Y(n13407) );
  nand2_1 U12729 ( .A(n13341), .B(n13297), .Y(n13100) );
  nor3_1 U12730 ( .A(n13367), .B(n13401), .C(n13369), .Y(n13297) );
  nor2_1 U12731 ( .A(n13227), .B(n13038), .Y(n13080) );
  inv_1 U12732 ( .A(n13180), .Y(n13038) );
  nor3_1 U12733 ( .A(n13408), .B(n13392), .C(n13380), .Y(n13180) );
  inv_1 U12734 ( .A(n13330), .Y(n13227) );
  nor2_1 U12735 ( .A(n13377), .B(n13409), .Y(n13330) );
  inv_1 U12736 ( .A(n13211), .Y(n13280) );
  nor2_1 U12737 ( .A(n13206), .B(n13391), .Y(n13211) );
  nand2_1 U12738 ( .A(n13397), .B(n13385), .Y(n13391) );
  inv_1 U12739 ( .A(n13337), .Y(n13206) );
  nor3_1 U12740 ( .A(n13408), .B(n13379), .C(n13380), .Y(n13337) );
  nand2_1 U12741 ( .A(n23979), .B(n13410), .Y(n13380) );
  a21oi_1 U12742 ( .A1(n13256), .A2(n13217), .B1(n13071), .Y(n13122) );
  inv_1 U12743 ( .A(n13305), .Y(n13071) );
  nand2_1 U12744 ( .A(n13259), .B(n13362), .Y(n13305) );
  nor2_1 U12745 ( .A(n13403), .B(n13378), .Y(n13362) );
  and4_1 U12746 ( .A(n13396), .B(n11751), .C(n24020), .D(n24003), .X(n13259)
         );
  nor2_1 U12747 ( .A(n13381), .B(n13378), .Y(n13217) );
  and2_0 U12748 ( .A(n13405), .B(n13400), .X(n13256) );
  nor3_1 U12749 ( .A(n24003), .B(n24020), .C(n11489), .Y(n13405) );
  nand4_1 U12750 ( .A(n13411), .B(n13412), .C(n13413), .D(n13414), .Y(n10409)
         );
  nor4_1 U12751 ( .A(n13415), .B(n13416), .C(n13417), .D(n13418), .Y(n13414)
         );
  a21oi_1 U12752 ( .A1(n13419), .A2(n13420), .B1(n12599), .Y(n13418) );
  nor4_1 U12753 ( .A(n13421), .B(n13422), .C(n13423), .D(n12603), .Y(n13420)
         );
  nand4_1 U12754 ( .A(n13424), .B(n13425), .C(n13426), .D(n13427), .Y(n13421)
         );
  nor4_1 U12755 ( .A(n13428), .B(n12610), .C(n13429), .D(n13430), .Y(n13419)
         );
  nand4_1 U12756 ( .A(n13431), .B(n12611), .C(n13432), .D(n13433), .Y(n13428)
         );
  and2_0 U12757 ( .A(n13434), .B(n13435), .X(n13417) );
  a21oi_1 U12758 ( .A1(n13436), .A2(n13437), .B1(n13438), .Y(n13416) );
  a221oi_1 U12759 ( .A1(n13439), .A2(n13440), .B1(n13441), .B2(n13442), .C1(
        n13443), .Y(n13413) );
  o22ai_1 U12760 ( .A1(n12596), .A2(n13444), .B1(n13445), .B2(n13446), .Y(
        n13443) );
  inv_1 U12761 ( .A(n13447), .Y(n13445) );
  inv_1 U12762 ( .A(n13448), .Y(n13440) );
  nor4_1 U12763 ( .A(n13449), .B(n12622), .C(n13450), .D(n13451), .Y(n13412)
         );
  nand4_1 U12764 ( .A(n13452), .B(n13453), .C(n13454), .D(n13455), .Y(n12622)
         );
  a222oi_1 U12765 ( .A1(n13456), .A2(n13434), .B1(n13457), .B2(n13458), .C1(
        n13459), .C2(n13460), .Y(n13455) );
  nand2_1 U12766 ( .A(n13461), .B(n12574), .Y(n13454) );
  nor2_1 U12767 ( .A(n12571), .B(n12620), .Y(n13449) );
  nor3_1 U12768 ( .A(n13462), .B(n13463), .C(n13464), .Y(n13411) );
  nand4_1 U12769 ( .A(n13465), .B(n13466), .C(n13467), .D(n13468), .Y(n10408)
         );
  nor3_1 U12770 ( .A(n13469), .B(n13470), .C(n13471), .Y(n13468) );
  o21ai_0 U12771 ( .A1(n13472), .A2(n13473), .B1(n13474), .Y(n13471) );
  o211ai_1 U12772 ( .A1(n13475), .A2(n13476), .B1(n13477), .C1(n13478), .Y(
        n13469) );
  o21ai_0 U12773 ( .A1(n13479), .A2(n13480), .B1(n12574), .Y(n13478) );
  nand4_1 U12774 ( .A(n13481), .B(n13482), .C(n13483), .D(n13484), .Y(n13480)
         );
  nor3_1 U12775 ( .A(n12609), .B(n13485), .C(n13430), .Y(n13484) );
  inv_1 U12776 ( .A(n12591), .Y(n13430) );
  nand4_1 U12777 ( .A(n13486), .B(n13487), .C(n13488), .D(n13489), .Y(n12609)
         );
  inv_1 U12778 ( .A(n13490), .Y(n13481) );
  nand4_1 U12779 ( .A(n12620), .B(n13491), .C(n12757), .D(n13492), .Y(n13479)
         );
  nor3_1 U12780 ( .A(n13493), .B(n13494), .C(n13495), .Y(n13492) );
  o21ai_0 U12781 ( .A1(n13496), .A2(n12602), .B1(n12617), .Y(n13477) );
  nor3_1 U12782 ( .A(n13497), .B(n13498), .C(n13499), .Y(n13467) );
  inv_1 U12783 ( .A(n13500), .Y(n13466) );
  or4_1 U12784 ( .A(n13501), .B(n13502), .C(n13503), .D(n13504), .X(n10407) );
  nand4_1 U12785 ( .A(n13505), .B(n13506), .C(n13507), .D(n13508), .Y(n13504)
         );
  a222oi_1 U12786 ( .A1(n13509), .A2(n12568), .B1(n13459), .B2(n13510), .C1(
        n13511), .C2(n13512), .Y(n13508) );
  inv_1 U12787 ( .A(n13491), .Y(n13459) );
  o21ai_0 U12788 ( .A1(n13513), .A2(n13514), .B1(n12574), .Y(n13507) );
  or4_1 U12789 ( .A(n12573), .B(n13493), .C(n13515), .D(n13516), .X(n13514) );
  nand4_1 U12790 ( .A(n13517), .B(n13518), .C(n13519), .D(n13520), .Y(n12573)
         );
  nor4_1 U12791 ( .A(n13521), .B(n13522), .C(n13523), .D(n13422), .Y(n13520)
         );
  nand4_1 U12792 ( .A(n13524), .B(n13525), .C(n13526), .D(n13527), .Y(n13521)
         );
  and3_1 U12793 ( .A(n13528), .B(n13529), .C(n13530), .X(n13519) );
  nor2_1 U12794 ( .A(n13531), .B(n13532), .Y(n13517) );
  nand4_1 U12795 ( .A(n13533), .B(n13476), .C(n13534), .D(n13535), .Y(n13513)
         );
  or3_1 U12796 ( .A(n13450), .B(n12575), .C(n13536), .X(n13503) );
  o22ai_1 U12797 ( .A1(n13537), .A2(n12757), .B1(n12599), .B2(n13538), .Y(
        n12575) );
  o22ai_1 U12798 ( .A1(n13537), .A2(n12613), .B1(n12571), .B2(n13539), .Y(
        n13450) );
  nand4_1 U12799 ( .A(n13540), .B(n12625), .C(n13541), .D(n13542), .Y(n10406)
         );
  nor4_1 U12800 ( .A(n13543), .B(n13544), .C(n13545), .D(n13546), .Y(n13542)
         );
  or3_1 U12801 ( .A(n13547), .B(n13548), .C(n13549), .X(n13543) );
  nor3_1 U12802 ( .A(n13550), .B(n13551), .C(n13552), .Y(n13541) );
  a21oi_1 U12803 ( .A1(n13553), .A2(n13554), .B1(n12596), .Y(n13552) );
  o22ai_1 U12804 ( .A1(n13555), .A2(n13556), .B1(n12599), .B2(n13557), .Y(
        n13550) );
  nor4_1 U12805 ( .A(n13558), .B(n13559), .C(n13560), .D(n13561), .Y(n13557)
         );
  nand4_1 U12806 ( .A(n13482), .B(n13562), .C(n12592), .D(n12606), .Y(n13561)
         );
  nand4_1 U12807 ( .A(n13563), .B(n13444), .C(n13564), .D(n13565), .Y(n13560)
         );
  nand4_1 U12808 ( .A(n13433), .B(n13529), .C(n13566), .D(n13567), .Y(n13559)
         );
  nand4_1 U12809 ( .A(n12757), .B(n13568), .C(n13569), .D(n13426), .Y(n13558)
         );
  nor2_1 U12810 ( .A(n13570), .B(n13571), .Y(n13569) );
  inv_1 U12811 ( .A(n13572), .Y(n13556) );
  a211oi_1 U12812 ( .A1(n13434), .A2(n13523), .B1(n13573), .C1(n13574), .Y(
        n12625) );
  a21oi_1 U12813 ( .A1(n13575), .A2(n13473), .B1(n13576), .Y(n13573) );
  a21oi_1 U12814 ( .A1(n13577), .A2(n13578), .B1(n12621), .Y(n13540) );
  nand4_1 U12815 ( .A(n13579), .B(n13474), .C(n13580), .D(n13581), .Y(n12621)
         );
  a22oi_1 U12816 ( .A1(n13495), .A2(n12568), .B1(n13515), .B2(n13582), .Y(
        n13580) );
  inv_1 U12817 ( .A(n13583), .Y(n13474) );
  o22ai_1 U12818 ( .A1(n13475), .A2(n13584), .B1(n13446), .B2(n13585), .Y(
        n13583) );
  inv_1 U12819 ( .A(n13586), .Y(n13579) );
  nand4_1 U12820 ( .A(n13587), .B(n12626), .C(n13588), .D(n13589), .Y(n10405)
         );
  nor4_1 U12821 ( .A(n13590), .B(n13591), .C(n13592), .D(n13593), .Y(n13589)
         );
  or3_1 U12822 ( .A(n13499), .B(n13594), .C(n13595), .X(n13590) );
  o211ai_1 U12823 ( .A1(n13596), .A2(n13597), .B1(n13598), .C1(n13599), .Y(
        n13499) );
  a21oi_1 U12824 ( .A1(n13441), .A2(n13442), .B1(n13551), .Y(n13599) );
  a221oi_1 U12825 ( .A1(n12601), .A2(n12619), .B1(n13600), .B2(n13458), .C1(
        n13601), .Y(n13588) );
  o22ai_1 U12826 ( .A1(n13448), .A2(n13602), .B1(n13603), .B2(n12599), .Y(
        n13601) );
  nor2_1 U12827 ( .A(n13604), .B(n13605), .Y(n13603) );
  nand4_1 U12828 ( .A(n13606), .B(n12592), .C(n13607), .D(n13608), .Y(n13605)
         );
  nor3_1 U12829 ( .A(n13609), .B(n13610), .C(n13515), .Y(n13608) );
  nand4_1 U12830 ( .A(n13611), .B(n13612), .C(n13476), .D(n13613), .Y(n13604)
         );
  nor4_1 U12831 ( .A(n13614), .B(n13511), .C(n13615), .D(n13522), .Y(n13613)
         );
  and4_1 U12832 ( .A(n13506), .B(n13616), .C(n13617), .D(n13618), .X(n12626)
         );
  a222oi_1 U12833 ( .A1(n13571), .A2(n12615), .B1(n13458), .B2(n13516), .C1(
        n13619), .C2(n13620), .Y(n13618) );
  inv_1 U12834 ( .A(n13621), .Y(n13516) );
  or2_0 U12835 ( .A(n13444), .B(n12596), .X(n13617) );
  a21oi_1 U12836 ( .A1(n12747), .A2(n13510), .B1(n13574), .Y(n13587) );
  or3_1 U12837 ( .A(n13622), .B(n13623), .C(n13624), .X(n13574) );
  and3_1 U12838 ( .A(n13625), .B(n13620), .C(n13626), .X(n13624) );
  nand4_1 U12839 ( .A(n13627), .B(n13628), .C(n13629), .D(n13630), .Y(n10404)
         );
  nor4_1 U12840 ( .A(n13631), .B(n13632), .C(n13633), .D(n13634), .Y(n13630)
         );
  nor2_1 U12841 ( .A(n12591), .B(n13635), .Y(n13634) );
  nor2_1 U12842 ( .A(n13636), .B(n13637), .Y(n12591) );
  a21oi_1 U12843 ( .A1(n13638), .A2(n13639), .B1(n12599), .Y(n13633) );
  nor4_1 U12844 ( .A(n13640), .B(n13641), .C(n13523), .D(n12601), .Y(n13639)
         );
  inv_1 U12845 ( .A(n13567), .Y(n12601) );
  nand3_1 U12846 ( .A(n13426), .B(n13642), .C(n13526), .Y(n13640) );
  nor4_1 U12847 ( .A(n13643), .B(n13644), .C(n13496), .D(n13645), .Y(n13638)
         );
  nand3_1 U12848 ( .A(n13533), .B(n13646), .C(n12611), .Y(n13643) );
  a21oi_1 U12849 ( .A1(n13647), .A2(n13529), .B1(n13648), .Y(n13632) );
  inv_1 U12850 ( .A(n13649), .Y(n13629) );
  o221ai_1 U12851 ( .A1(n13650), .A2(n13555), .B1(n12593), .B2(n13483), .C1(
        n12624), .Y(n13649) );
  a221oi_1 U12852 ( .A1(n13651), .A2(n13578), .B1(n13652), .B2(n13653), .C1(
        n13654), .Y(n12624) );
  o211ai_1 U12853 ( .A1(n13448), .A2(n13597), .B1(n13655), .C1(n13505), .Y(
        n13654) );
  inv_1 U12854 ( .A(n13476), .Y(n13651) );
  nor3_1 U12855 ( .A(n13536), .B(n13451), .C(n13656), .Y(n13628) );
  o221ai_1 U12856 ( .A1(n13438), .A2(n13562), .B1(n13635), .B2(n13657), .C1(
        n13658), .Y(n13451) );
  a21oi_1 U12857 ( .A1(n13659), .A2(n13512), .B1(n13660), .Y(n13658) );
  inv_1 U12858 ( .A(n13473), .Y(n13659) );
  o21ai_0 U12859 ( .A1(n13446), .A2(n12605), .B1(n13661), .Y(n13536) );
  inv_1 U12860 ( .A(n13662), .Y(n13661) );
  nor3_1 U12861 ( .A(n13663), .B(n13544), .C(n13664), .Y(n13627) );
  o211ai_1 U12862 ( .A1(n13537), .A2(n13491), .B1(n13665), .C1(n13666), .Y(
        n13544) );
  a222oi_1 U12863 ( .A1(n13667), .A2(n12574), .B1(n13461), .B2(n13439), .C1(
        n12616), .C2(n13582), .Y(n13666) );
  nand4_1 U12864 ( .A(n13668), .B(n13669), .C(n13670), .D(n13671), .Y(n10403)
         );
  a221oi_1 U12865 ( .A1(n13447), .A2(n13672), .B1(n13461), .B2(n13439), .C1(
        n13673), .Y(n13671) );
  o21ai_0 U12866 ( .A1(n12599), .A2(n13674), .B1(n13675), .Y(n13673) );
  nor4_1 U12867 ( .A(n13676), .B(n13677), .C(n13678), .D(n13572), .Y(n13674)
         );
  nand2_1 U12868 ( .A(n12611), .B(n13679), .Y(n13572) );
  nand3_1 U12869 ( .A(n13483), .B(n13437), .C(n13680), .Y(n13677) );
  inv_1 U12870 ( .A(n13681), .Y(n13680) );
  nand4_1 U12871 ( .A(n13553), .B(n13488), .C(n13562), .D(n13682), .Y(n13676)
         );
  and3_1 U12872 ( .A(n13444), .B(n13527), .C(n13538), .X(n13682) );
  inv_1 U12873 ( .A(n13683), .Y(n13461) );
  nand3_1 U12874 ( .A(n13476), .B(n13530), .C(n13584), .Y(n13447) );
  a222oi_1 U12875 ( .A1(n13684), .A2(n13442), .B1(n12616), .B2(n12617), .C1(
        n13685), .C2(n13510), .Y(n13670) );
  inv_1 U12876 ( .A(n12613), .Y(n13685) );
  nor3_1 U12877 ( .A(n13500), .B(n13686), .C(n13497), .Y(n13669) );
  or4_1 U12878 ( .A(n13687), .B(n13656), .C(n13688), .D(n13547), .X(n13497) );
  o22ai_1 U12879 ( .A1(n13635), .A2(n13533), .B1(n13555), .B2(n13621), .Y(
        n13547) );
  o21ai_0 U12880 ( .A1(n13563), .A2(n13689), .B1(n13690), .Y(n13688) );
  inv_1 U12881 ( .A(n13691), .Y(n13690) );
  o21ai_0 U12882 ( .A1(n12596), .A2(n12606), .B1(n13692), .Y(n13656) );
  nand4_1 U12883 ( .A(n13693), .B(n13694), .C(n13695), .D(n13696), .Y(n13500)
         );
  a221oi_1 U12884 ( .A1(n13697), .A2(n13434), .B1(n13571), .B2(n12619), .C1(
        n13662), .Y(n13696) );
  o22ai_1 U12885 ( .A1(n12571), .A2(n13698), .B1(n13472), .B2(n13699), .Y(
        n13662) );
  o21ai_0 U12886 ( .A1(n13511), .A2(n13653), .B1(n13512), .Y(n13695) );
  nor3_1 U12887 ( .A(n13700), .B(n13546), .C(n13701), .Y(n13668) );
  o221ai_1 U12888 ( .A1(n13537), .A2(n12595), .B1(n13597), .B2(n13486), .C1(
        n13702), .Y(n13546) );
  nand2_1 U12889 ( .A(n13636), .B(n12568), .Y(n13702) );
  nand4_1 U12890 ( .A(n13703), .B(n13704), .C(n13705), .D(n13706), .Y(n10402)
         );
  nor4_1 U12891 ( .A(n13707), .B(n13708), .C(n13709), .D(n13710), .Y(n13706)
         );
  a21oi_1 U12892 ( .A1(n13612), .A2(n13699), .B1(n13576), .Y(n13710) );
  a21oi_1 U12893 ( .A1(n13711), .A2(n13712), .B1(n12599), .Y(n13708) );
  nor4_1 U12894 ( .A(n13713), .B(n13637), .C(n12602), .D(n13511), .Y(n13712)
         );
  inv_1 U12895 ( .A(n13714), .Y(n13637) );
  nand3_1 U12896 ( .A(n13527), .B(n13491), .C(n13528), .Y(n13713) );
  nor4_1 U12897 ( .A(n13715), .B(n13716), .C(n13717), .D(n13490), .Y(n13711)
         );
  nand3_1 U12898 ( .A(n13606), .B(n13718), .C(n13719), .Y(n13490) );
  inv_1 U12899 ( .A(n13645), .Y(n13719) );
  nand4_1 U12900 ( .A(n13431), .B(n13553), .C(n12595), .D(n13444), .Y(n13645)
         );
  nand3_1 U12901 ( .A(n13720), .B(n13721), .C(n13722), .Y(n13444) );
  and4_1 U12902 ( .A(n12604), .B(n13433), .C(n13683), .D(n13723), .X(n13606)
         );
  nand3_1 U12903 ( .A(n13724), .B(n13721), .C(n13725), .Y(n13683) );
  nand3_1 U12904 ( .A(n13533), .B(n13538), .C(n13473), .Y(n13715) );
  o22ai_1 U12905 ( .A1(n13537), .A2(n13726), .B1(n13648), .B2(n13567), .Y(
        n13707) );
  a221oi_1 U12906 ( .A1(n13684), .A2(n13458), .B1(n13609), .B2(n13434), .C1(
        n13727), .Y(n13705) );
  o22ai_1 U12907 ( .A1(n13483), .A2(n12593), .B1(n13555), .B2(n13728), .Y(
        n13727) );
  inv_1 U12908 ( .A(n13489), .Y(n13609) );
  nor4_1 U12909 ( .A(n13586), .B(n12623), .C(n13687), .D(n13729), .Y(n13704)
         );
  inv_1 U12910 ( .A(n13465), .Y(n13729) );
  nor4_1 U12911 ( .A(n13730), .B(n13594), .C(n13731), .D(n13732), .Y(n13465)
         );
  or4_1 U12912 ( .A(n13733), .B(n13734), .C(n13735), .D(n13622), .X(n13732) );
  inv_1 U12913 ( .A(n13453), .Y(n13735) );
  a21oi_1 U12914 ( .A1(n13650), .A2(n13679), .B1(n13555), .Y(n13734) );
  o22ai_1 U12915 ( .A1(n13597), .A2(n13448), .B1(n12596), .B2(n13736), .Y(
        n13733) );
  inv_1 U12916 ( .A(n13737), .Y(n13731) );
  a21oi_1 U12917 ( .A1(n13738), .A2(n12619), .B1(n13660), .Y(n13737) );
  o21ai_0 U12918 ( .A1(n12572), .A2(n13648), .B1(n13739), .Y(n13660) );
  nand3_1 U12919 ( .A(n13725), .B(n13724), .C(n13740), .Y(n12572) );
  o221ai_1 U12920 ( .A1(n12596), .A2(n12613), .B1(n13555), .B2(n12611), .C1(
        n13452), .Y(n13594) );
  nand4_1 U12921 ( .A(n13741), .B(n13742), .C(n13620), .D(n13743), .Y(n13452)
         );
  nand4_1 U12922 ( .A(n13744), .B(n13745), .C(n13746), .D(n13747), .Y(n13687)
         );
  nor3_1 U12923 ( .A(n13748), .B(n13749), .C(n13750), .Y(n13747) );
  inv_1 U12924 ( .A(n13665), .Y(n13750) );
  nor2_1 U12925 ( .A(n13415), .B(n13751), .Y(n13665) );
  and4_1 U12926 ( .A(n13752), .B(n13741), .C(n13439), .D(n13740), .X(n13751)
         );
  inv_1 U12927 ( .A(n13753), .Y(n13415) );
  o22ai_1 U12928 ( .A1(n13635), .A2(n13564), .B1(n13438), .B2(n13754), .Y(
        n13748) );
  nor3_1 U12929 ( .A(n13623), .B(n13631), .C(n13755), .Y(n13746) );
  o221ai_1 U12930 ( .A1(n13756), .A2(n13566), .B1(n12599), .B2(n13563), .C1(
        n13757), .Y(n12623) );
  nand2_1 U12931 ( .A(n13577), .B(n13672), .Y(n13757) );
  o221ai_1 U12932 ( .A1(n12596), .A2(n13524), .B1(n13602), .B2(n13646), .C1(
        n13758), .Y(n13586) );
  nor4_1 U12933 ( .A(n13759), .B(n13545), .C(n13592), .D(n13701), .Y(n13703)
         );
  o22ai_1 U12934 ( .A1(n13576), .A2(n13525), .B1(n13635), .B2(n13760), .Y(
        n13701) );
  o22ai_1 U12935 ( .A1(n13602), .A2(n13486), .B1(n13761), .B2(n12593), .Y(
        n13592) );
  nor2_1 U12936 ( .A(n13636), .B(n13495), .Y(n13761) );
  inv_1 U12937 ( .A(n13657), .Y(n13495) );
  nor3_1 U12938 ( .A(n13762), .B(n13763), .C(n13764), .Y(n13636) );
  inv_1 U12939 ( .A(n13765), .Y(n13545) );
  a221oi_1 U12940 ( .A1(n13582), .A2(n13766), .B1(n12617), .B2(n13641), .C1(
        n13767), .Y(n13765) );
  o221ai_1 U12941 ( .A1(n13488), .A2(n13446), .B1(n13768), .B2(n12599), .C1(
        n13769), .Y(n13767) );
  inv_1 U12942 ( .A(n13770), .Y(n13759) );
  nand4_1 U12943 ( .A(n13771), .B(n13772), .C(n13773), .D(n13774), .Y(n10401)
         );
  nor3_1 U12944 ( .A(n13775), .B(n13755), .C(n13776), .Y(n13774) );
  a21oi_1 U12945 ( .A1(n13777), .A2(n13778), .B1(n12599), .Y(n13776) );
  nor4_1 U12946 ( .A(n12747), .B(n13641), .C(n13779), .D(n13457), .Y(n13778)
         );
  inv_1 U12947 ( .A(n13679), .Y(n13457) );
  nor4_1 U12948 ( .A(n13684), .B(n13531), .C(n13780), .D(n13681), .Y(n13777)
         );
  nand4_1 U12949 ( .A(n13482), .B(n13718), .C(n13647), .D(n13657), .Y(n13681)
         );
  nor3_1 U12950 ( .A(n13600), .B(n13614), .C(n12610), .Y(n13482) );
  inv_1 U12951 ( .A(n13607), .Y(n13780) );
  nor4_1 U12952 ( .A(n12608), .B(n13494), .C(n13523), .D(n13766), .Y(n13607)
         );
  inv_1 U12953 ( .A(n13781), .Y(n13523) );
  nand3_1 U12954 ( .A(n13529), .B(n13527), .C(n13650), .Y(n12608) );
  nand2_1 U12955 ( .A(n13782), .B(n13783), .Y(n13527) );
  nand3_1 U12956 ( .A(n13784), .B(n13785), .C(n13786), .Y(n13529) );
  nand4_1 U12957 ( .A(n13567), .B(n13612), .C(n13566), .D(n13787), .Y(n13531)
         );
  nor3_1 U12958 ( .A(n12603), .B(n13788), .C(n13615), .Y(n13787) );
  inv_1 U12959 ( .A(n13575), .Y(n13615) );
  inv_1 U12960 ( .A(n13789), .Y(n13684) );
  a21oi_1 U12961 ( .A1(n12620), .A2(n13433), .B1(n12571), .Y(n13775) );
  a222oi_1 U12962 ( .A1(n13423), .A2(n13460), .B1(n13610), .B2(n12568), .C1(
        n13511), .C2(n13652), .Y(n13773) );
  inv_1 U12963 ( .A(n13426), .Y(n13511) );
  inv_1 U12964 ( .A(n13524), .Y(n13423) );
  nor3_1 U12965 ( .A(n13593), .B(n13730), .C(n13691), .Y(n13772) );
  o21ai_0 U12966 ( .A1(n13689), .A2(n13436), .B1(n13790), .Y(n13691) );
  o21ai_0 U12967 ( .A1(n13689), .A2(n13424), .B1(n13791), .Y(n13730) );
  nand4_1 U12968 ( .A(n13693), .B(n13655), .C(n13792), .D(n13793), .Y(n13593)
         );
  a22oi_1 U12969 ( .A1(n13577), .A2(n13672), .B1(n13697), .B2(n13439), .Y(
        n13793) );
  inv_1 U12970 ( .A(n13530), .Y(n13577) );
  nand2_1 U12971 ( .A(n13794), .B(n13785), .Y(n13530) );
  o21ai_0 U12972 ( .A1(n12616), .A2(n13485), .B1(n12574), .Y(n13792) );
  inv_1 U12973 ( .A(n13528), .Y(n12616) );
  nand2_1 U12974 ( .A(n13795), .B(n13794), .Y(n13528) );
  inv_1 U12975 ( .A(n13796), .Y(n13655) );
  a21oi_1 U12976 ( .A1(n13538), .A2(n13525), .B1(n13576), .Y(n13796) );
  nor3_1 U12977 ( .A(n13797), .B(n13591), .C(n13664), .Y(n13771) );
  or4_1 U12978 ( .A(n13798), .B(n13799), .C(n13800), .D(n13801), .X(n13664) );
  o221ai_1 U12979 ( .A1(n13602), .A2(n13596), .B1(n13611), .B2(n13648), .C1(
        n13581), .Y(n13801) );
  a21oi_1 U12980 ( .A1(n12617), .A2(n13522), .B1(n13802), .Y(n13581) );
  nor2_1 U12981 ( .A(n13760), .B(n12593), .Y(n13800) );
  a21oi_1 U12982 ( .A1(n13486), .A2(n13489), .B1(n13597), .Y(n13798) );
  or3_1 U12983 ( .A(n13803), .B(n13804), .C(n13805), .X(n13591) );
  inv_1 U12984 ( .A(n13806), .Y(n13805) );
  a222oi_1 U12985 ( .A1(n12602), .A2(n12617), .B1(n13738), .B2(n12615), .C1(
        n13496), .C2(n13582), .Y(n13806) );
  inv_1 U12986 ( .A(n13437), .Y(n13496) );
  inv_1 U12987 ( .A(n13642), .Y(n12602) );
  nand4_1 U12988 ( .A(n13807), .B(n13808), .C(n13809), .D(n13810), .Y(n10400)
         );
  nor4_1 U12989 ( .A(n13755), .B(n13551), .C(n13799), .D(n13622), .Y(n13810)
         );
  nor2_1 U12990 ( .A(n13427), .B(n13756), .Y(n13622) );
  nor2_1 U12991 ( .A(n13736), .B(n13537), .Y(n13799) );
  a21oi_1 U12992 ( .A1(n13728), .A2(n13789), .B1(n13555), .Y(n13551) );
  inv_1 U12993 ( .A(n13442), .Y(n13555) );
  and2_0 U12994 ( .A(n13570), .B(n12617), .X(n13755) );
  a221oi_1 U12995 ( .A1(n13811), .A2(n13460), .B1(n13620), .B2(n13812), .C1(
        n13813), .Y(n13809) );
  o22ai_1 U12996 ( .A1(n13648), .A2(n13567), .B1(n12599), .B2(n13814), .Y(
        n13813) );
  nor4_1 U12997 ( .A(n13815), .B(n13816), .C(n13644), .D(n13435), .Y(n13814)
         );
  o21ai_0 U12998 ( .A1(n13817), .A2(n13818), .B1(n13486), .Y(n13435) );
  nand4_1 U12999 ( .A(n13819), .B(n13725), .C(n13820), .D(n13821), .Y(n13486)
         );
  nand4_1 U13000 ( .A(n13563), .B(n13621), .C(n13822), .D(n13823), .Y(n13644)
         );
  nor4_1 U13001 ( .A(n13824), .B(n13738), .C(n12610), .D(n13716), .Y(n13823)
         );
  nand2_1 U13002 ( .A(n12757), .B(n13584), .Y(n13716) );
  o32ai_1 U13003 ( .A1(n13825), .A2(n13826), .A3(n13827), .B1(n13828), .B2(
        n13829), .Y(n12610) );
  nand2_1 U13004 ( .A(n13743), .B(n13830), .Y(n13829) );
  inv_1 U13005 ( .A(n13539), .Y(n13738) );
  nand3_1 U13006 ( .A(n13831), .B(n13832), .C(n13833), .Y(n13539) );
  inv_1 U13007 ( .A(n13488), .Y(n13824) );
  nor3_1 U13008 ( .A(n13494), .B(n13571), .C(n13441), .Y(n13822) );
  inv_1 U13009 ( .A(n13566), .Y(n13441) );
  nand3_1 U13010 ( .A(n13786), .B(n13785), .C(n13834), .Y(n13566) );
  inv_1 U13011 ( .A(n13534), .Y(n13571) );
  inv_1 U13012 ( .A(n13432), .Y(n13494) );
  nand3_1 U13013 ( .A(n13835), .B(n13833), .C(n13836), .Y(n13621) );
  nand3_1 U13014 ( .A(n13518), .B(n12613), .C(n13718), .Y(n13816) );
  and2_0 U13015 ( .A(n13554), .B(n13568), .X(n13718) );
  nand3_1 U13016 ( .A(n13837), .B(n13832), .C(n13838), .Y(n12613) );
  nor4_1 U13017 ( .A(n12618), .B(n13839), .C(n13779), .D(n13641), .Y(n13518)
         );
  inv_1 U13018 ( .A(n13760), .Y(n13839) );
  inv_1 U13019 ( .A(n13433), .Y(n12618) );
  nand2_1 U13020 ( .A(n13784), .B(n13783), .Y(n13433) );
  nand4_1 U13021 ( .A(n13657), .B(n13436), .C(n13679), .D(n13840), .Y(n13815)
         );
  and3_1 U13022 ( .A(n13448), .B(n13424), .C(n13476), .X(n13840) );
  nand3_1 U13023 ( .A(n13838), .B(n13837), .C(n13841), .Y(n13424) );
  nand3_1 U13024 ( .A(n13833), .B(n13831), .C(n13841), .Y(n13448) );
  nand4_1 U13025 ( .A(n13842), .B(n13843), .C(n13844), .D(n13845), .Y(n13679)
         );
  nand3_1 U13026 ( .A(n13846), .B(n13847), .C(n13795), .Y(n13567) );
  nand3_1 U13027 ( .A(n13533), .B(n13535), .C(n12604), .Y(n13812) );
  nand2_1 U13028 ( .A(n12606), .B(n12595), .Y(n13811) );
  nand3_1 U13029 ( .A(n13848), .B(n13740), .C(n13720), .Y(n12595) );
  a221oi_1 U13030 ( .A1(n13600), .A2(n13458), .B1(n13766), .B2(n12617), .C1(
        n13849), .Y(n13808) );
  o22ai_1 U13031 ( .A1(n13597), .A2(n13425), .B1(n13472), .B2(n13538), .Y(
        n13849) );
  nand3_1 U13032 ( .A(n13850), .B(n13847), .C(n13846), .Y(n13538) );
  inv_1 U13033 ( .A(n13434), .Y(n13597) );
  inv_1 U13034 ( .A(n13526), .Y(n13766) );
  nor3_1 U13035 ( .A(n13803), .B(n13463), .C(n13501), .Y(n13807) );
  nand4_1 U13036 ( .A(n13739), .B(n13675), .C(n13851), .D(n13852), .Y(n13501)
         );
  a211oi_1 U13037 ( .A1(n13853), .A2(n13510), .B1(n13854), .C1(n13549), .Y(
        n13852) );
  o221ai_1 U13038 ( .A1(n13689), .A2(n13437), .B1(n12596), .B2(n13726), .C1(
        n13693), .Y(n13549) );
  nand2_1 U13039 ( .A(n13855), .B(n13856), .Y(n13693) );
  o32ai_1 U13040 ( .A1(n13576), .A2(n13826), .A3(n13763), .B1(n13857), .B2(
        n13858), .Y(n13856) );
  inv_1 U13041 ( .A(n13830), .Y(n13857) );
  nand3_1 U13042 ( .A(n13833), .B(n13832), .C(n13859), .Y(n13437) );
  o22ai_1 U13043 ( .A1(n13635), .A2(n13714), .B1(n13756), .B2(n12611), .Y(
        n13854) );
  nand3_1 U13044 ( .A(n13860), .B(n13841), .C(n13842), .Y(n12611) );
  inv_1 U13045 ( .A(n13861), .Y(n13851) );
  o21ai_0 U13046 ( .A1(n13431), .A2(n13446), .B1(n13744), .Y(n13861) );
  nand3_1 U13047 ( .A(n13862), .B(n13725), .C(n13742), .Y(n13431) );
  nand4_1 U13048 ( .A(n13505), .B(n13791), .C(n13863), .D(n13864), .Y(n13463)
         );
  nor3_1 U13049 ( .A(n13865), .B(n13548), .C(n13498), .Y(n13864) );
  o221ai_1 U13050 ( .A1(n12571), .A2(n13611), .B1(n13576), .B2(n13575), .C1(
        n13866), .Y(n13498) );
  nand2_1 U13051 ( .A(n13667), .B(n13512), .Y(n13866) );
  inv_1 U13052 ( .A(n13612), .Y(n13667) );
  nand3_1 U13053 ( .A(n13867), .B(n13868), .C(n13794), .Y(n13612) );
  and2_0 U13054 ( .A(n13834), .B(n13869), .X(n13794) );
  o22ai_1 U13055 ( .A1(n13438), .A2(n13642), .B1(n13602), .B2(n12612), .Y(
        n13548) );
  o22ai_1 U13056 ( .A1(n13648), .A2(n13768), .B1(n13756), .B2(n13650), .Y(
        n13865) );
  nand2_1 U13057 ( .A(n13870), .B(n13841), .Y(n13650) );
  a21oi_1 U13058 ( .A1(n13522), .A2(n13582), .B1(n13802), .Y(n13863) );
  inv_1 U13059 ( .A(n13694), .Y(n13802) );
  o21ai_0 U13060 ( .A1(n13871), .A2(n13872), .B1(n13725), .Y(n13694) );
  nor3_1 U13061 ( .A(n13873), .B(n13874), .C(n13648), .Y(n13872) );
  nor3_1 U13062 ( .A(n13825), .B(n13537), .C(n13764), .Y(n13871) );
  inv_1 U13063 ( .A(n13754), .Y(n13522) );
  nand3_1 U13064 ( .A(n13782), .B(n13850), .C(n13869), .Y(n13754) );
  nand4_1 U13065 ( .A(n13855), .B(n12615), .C(n13721), .D(n13830), .Y(n13791)
         );
  nand2_1 U13066 ( .A(n13620), .B(n13610), .Y(n13505) );
  inv_1 U13067 ( .A(n13564), .Y(n13610) );
  nand4_1 U13068 ( .A(n13875), .B(n13758), .C(n13745), .D(n13876), .Y(n13803)
         );
  a22oi_1 U13069 ( .A1(n13422), .A2(n13578), .B1(n13653), .B2(n13512), .Y(
        n13876) );
  inv_1 U13070 ( .A(n13585), .Y(n13422) );
  nand3_1 U13071 ( .A(n12615), .B(n13838), .C(n13877), .Y(n13758) );
  nand4_1 U13072 ( .A(n13878), .B(n13879), .C(n13880), .D(n13881), .Y(n10399)
         );
  nor3_1 U13073 ( .A(n13882), .B(n13709), .C(n13883), .Y(n13881) );
  a21oi_1 U13074 ( .A1(n13760), .A2(n13657), .B1(n12593), .Y(n13883) );
  nand3_1 U13075 ( .A(n13721), .B(n13830), .C(n13884), .Y(n13657) );
  nand4_1 U13076 ( .A(n13834), .B(n13850), .C(n13885), .D(n13886), .Y(n13760)
         );
  inv_1 U13077 ( .A(n13875), .Y(n13709) );
  nand2_1 U13078 ( .A(n13493), .B(n12617), .Y(n13875) );
  inv_1 U13079 ( .A(n13562), .Y(n13493) );
  nand3_1 U13080 ( .A(n13848), .B(n13740), .C(n13884), .Y(n13562) );
  o22ai_1 U13081 ( .A1(n12599), .A2(n13887), .B1(n13475), .B2(n13585), .Y(
        n13882) );
  nand2_1 U13082 ( .A(n13888), .B(n13782), .Y(n13585) );
  nor4_1 U13083 ( .A(n13889), .B(n13890), .C(n13619), .D(n13515), .Y(n13887)
         );
  inv_1 U13084 ( .A(n13436), .Y(n13515) );
  nand2_1 U13085 ( .A(n13877), .B(n13835), .Y(n13436) );
  inv_1 U13086 ( .A(n13533), .Y(n13619) );
  nand2_1 U13087 ( .A(n13870), .B(n13891), .Y(n13533) );
  nand3_1 U13088 ( .A(n13699), .B(n13426), .C(n13564), .Y(n13890) );
  nand2_1 U13089 ( .A(n13892), .B(n13843), .Y(n13564) );
  nand2_1 U13090 ( .A(n13893), .B(n13831), .Y(n13426) );
  nand3_1 U13091 ( .A(n13836), .B(n13860), .C(n13859), .Y(n13699) );
  or4_1 U13092 ( .A(n13894), .B(n13678), .C(n13532), .D(n13697), .X(n13889) );
  inv_1 U13093 ( .A(n12612), .Y(n13697) );
  nand3_1 U13094 ( .A(n13836), .B(n13831), .C(n13895), .Y(n12612) );
  nand3_1 U13095 ( .A(n13611), .B(n13432), .C(n13596), .Y(n13532) );
  inv_1 U13096 ( .A(n13896), .Y(n13596) );
  o21ai_0 U13097 ( .A1(n13817), .A2(n13818), .B1(n13425), .Y(n13896) );
  nand3_1 U13098 ( .A(n13834), .B(n13786), .C(n13795), .Y(n13425) );
  nand3_1 U13099 ( .A(n13869), .B(n13782), .C(n13795), .Y(n13432) );
  nand2_1 U13100 ( .A(n13888), .B(n13846), .Y(n13611) );
  nand4_1 U13101 ( .A(n13491), .B(n13714), .C(n12620), .D(n13897), .Y(n13678)
         );
  and2_0 U13102 ( .A(n13487), .B(n13726), .X(n13897) );
  inv_1 U13103 ( .A(n13485), .Y(n13726) );
  nor3_1 U13104 ( .A(n13898), .B(n13826), .C(n13825), .Y(n13485) );
  inv_1 U13105 ( .A(n13724), .Y(n13826) );
  nand3_1 U13106 ( .A(n13743), .B(n13830), .C(n13740), .Y(n13487) );
  nand4_1 U13107 ( .A(n13752), .B(n13830), .C(n13820), .D(n13821), .Y(n12620)
         );
  nand3_1 U13108 ( .A(n13742), .B(n13884), .C(n13741), .Y(n13714) );
  nand3_1 U13109 ( .A(n13720), .B(n13721), .C(n13819), .Y(n13491) );
  inv_1 U13110 ( .A(n13698), .Y(n13894) );
  a21oi_1 U13111 ( .A1(n13838), .A2(n13877), .B1(n13899), .Y(n13698) );
  inv_1 U13112 ( .A(n13768), .Y(n13899) );
  nand3_1 U13113 ( .A(n13837), .B(n13831), .C(n13836), .Y(n13768) );
  and3_1 U13114 ( .A(n13844), .B(n13845), .C(n13836), .X(n13877) );
  a221oi_1 U13115 ( .A1(n13614), .A2(n12568), .B1(n12603), .B2(n13458), .C1(
        n13900), .Y(n13880) );
  o22ai_1 U13116 ( .A1(n13648), .A2(n13534), .B1(n13781), .B2(n13602), .Y(
        n13900) );
  nand2_1 U13117 ( .A(n13834), .B(n13888), .Y(n13781) );
  and3_1 U13118 ( .A(n13885), .B(n13886), .C(n13785), .X(n13888) );
  nand2_1 U13119 ( .A(n13859), .B(n13893), .Y(n13534) );
  inv_1 U13120 ( .A(n13728), .Y(n12603) );
  nand2_1 U13121 ( .A(n13901), .B(n13786), .Y(n13728) );
  inv_1 U13122 ( .A(n13535), .Y(n13614) );
  nand4_1 U13123 ( .A(n13819), .B(n13720), .C(n13820), .D(n13821), .Y(n13535)
         );
  nor4_1 U13124 ( .A(n13902), .B(n13464), .C(n13462), .D(n13502), .Y(n13879)
         );
  nand4_1 U13125 ( .A(n13770), .B(n13692), .C(n13903), .D(n13904), .Y(n13502)
         );
  nor3_1 U13126 ( .A(n13905), .B(n13631), .C(n13906), .Y(n13904) );
  inv_1 U13127 ( .A(n13745), .Y(n13906) );
  nand4_1 U13128 ( .A(n13439), .B(n13626), .C(n13724), .D(n13743), .Y(n13745)
         );
  nor4_1 U13129 ( .A(n13907), .B(n13828), .C(n13602), .D(n13762), .Y(n13631)
         );
  o22ai_1 U13130 ( .A1(n13576), .A2(n13473), .B1(n13438), .B2(n13642), .Y(
        n13905) );
  nand2_1 U13131 ( .A(n13893), .B(n13842), .Y(n13642) );
  nand2_1 U13132 ( .A(n13841), .B(n13892), .Y(n13473) );
  inv_1 U13133 ( .A(n13595), .Y(n13903) );
  o221ai_1 U13134 ( .A1(n13537), .A2(n13554), .B1(n13438), .B2(n13563), .C1(
        n13753), .Y(n13595) );
  nand4_1 U13135 ( .A(n13752), .B(n13439), .C(n13626), .D(n13862), .Y(n13753)
         );
  nand3_1 U13136 ( .A(n13891), .B(n13838), .C(n13895), .Y(n13563) );
  nand3_1 U13137 ( .A(n13848), .B(n13725), .C(n13742), .Y(n13554) );
  and2_0 U13138 ( .A(n13769), .B(n13908), .X(n13692) );
  nand4_1 U13139 ( .A(n13752), .B(n13626), .C(n13722), .D(n13578), .Y(n13908)
         );
  inv_1 U13140 ( .A(n13446), .Y(n13578) );
  nand4_1 U13141 ( .A(n13819), .B(n12615), .C(n13740), .D(n13743), .Y(n13769)
         );
  inv_1 U13142 ( .A(n13907), .Y(n13819) );
  a22oi_1 U13143 ( .A1(n13442), .A2(n13600), .B1(n13652), .B2(n13653), .Y(
        n13770) );
  inv_1 U13144 ( .A(n13565), .Y(n13653) );
  nand2_1 U13145 ( .A(n13909), .B(n13841), .Y(n13565) );
  inv_1 U13146 ( .A(n13576), .Y(n13652) );
  nand2_1 U13147 ( .A(n13910), .B(n13911), .Y(n13576) );
  and3_1 U13148 ( .A(n13741), .B(n13626), .C(n13752), .X(n13600) );
  nand4_1 U13149 ( .A(n13912), .B(n13913), .C(n13914), .D(n13598), .Y(n13462)
         );
  a22oi_1 U13150 ( .A1(n13582), .A2(n13641), .B1(n13434), .B2(n13779), .Y(
        n13598) );
  inv_1 U13151 ( .A(n13646), .Y(n13779) );
  nand3_1 U13152 ( .A(n13786), .B(n13846), .C(n13795), .Y(n13646) );
  and2_0 U13153 ( .A(n13915), .B(n13916), .X(n13795) );
  o21ai_0 U13154 ( .A1(n13917), .A2(n12599), .B1(n13918), .Y(n13434) );
  and2_0 U13155 ( .A(n13901), .B(n13869), .X(n13641) );
  and3_1 U13156 ( .A(n13867), .B(n13868), .C(n13784), .X(n13901) );
  a21oi_1 U13157 ( .A1(n13919), .A2(n13512), .B1(n13749), .Y(n13914) );
  o21ai_0 U13158 ( .A1(n13475), .A2(n12605), .B1(n13616), .Y(n13749) );
  nand4_1 U13159 ( .A(n13920), .B(n13510), .C(n13921), .D(n13922), .Y(n13616)
         );
  nand2_1 U13160 ( .A(n13909), .B(n13891), .Y(n12605) );
  inv_1 U13161 ( .A(n13525), .Y(n13919) );
  nand3_1 U13162 ( .A(n13869), .B(n13850), .C(n13784), .Y(n13525) );
  and2_0 U13163 ( .A(n13923), .B(n13844), .X(n13784) );
  and2_0 U13164 ( .A(n13885), .B(n13924), .X(n13869) );
  inv_1 U13165 ( .A(n13686), .Y(n13913) );
  o22ai_1 U13166 ( .A1(n13602), .A2(n13489), .B1(n13635), .B2(n12604), .Y(
        n13686) );
  nand2_1 U13167 ( .A(n13625), .B(n13740), .Y(n12604) );
  nand3_1 U13168 ( .A(n13855), .B(n13721), .C(n13741), .Y(n13489) );
  inv_1 U13169 ( .A(n13470), .Y(n13912) );
  o22ai_1 U13170 ( .A1(n13689), .A2(n13526), .B1(n12571), .B2(n13647), .Y(
        n13470) );
  nand3_1 U13171 ( .A(n13860), .B(n13891), .C(n13842), .Y(n13647) );
  inv_1 U13172 ( .A(n12619), .Y(n12571) );
  o21ai_0 U13173 ( .A1(n13917), .A2(n12599), .B1(n13925), .Y(n12619) );
  nand3_1 U13174 ( .A(n13782), .B(n13847), .C(n13785), .Y(n13526) );
  and2_0 U13175 ( .A(n13926), .B(n13927), .X(n13785) );
  nor3_1 U13176 ( .A(n13928), .B(n13929), .C(n13930), .Y(n13847) );
  and2_0 U13177 ( .A(n13923), .B(n13931), .X(n13782) );
  nor3_1 U13178 ( .A(n10624), .B(n24008), .C(n12968), .Y(n13923) );
  inv_1 U13179 ( .A(n12617), .Y(n13689) );
  o21ai_0 U13180 ( .A1(n13910), .A2(n12599), .B1(n13918), .Y(n12617) );
  o221ai_1 U13181 ( .A1(n13537), .A2(n13553), .B1(n13475), .B2(n13488), .C1(
        n13932), .Y(n13464) );
  inv_1 U13182 ( .A(n13933), .Y(n13932) );
  o211ai_1 U13183 ( .A1(n13568), .A2(n13635), .B1(n13790), .C1(n13506), .Y(
        n13933) );
  nand2_1 U13184 ( .A(n13570), .B(n13582), .Y(n13506) );
  and3_1 U13185 ( .A(n13860), .B(n13843), .C(n13842), .X(n13570) );
  inv_1 U13186 ( .A(n13934), .Y(n13842) );
  nand4_1 U13187 ( .A(n13752), .B(n13722), .C(n13582), .D(n13740), .Y(n13790)
         );
  inv_1 U13188 ( .A(n13763), .Y(n13740) );
  nand2_1 U13189 ( .A(n13935), .B(n13821), .Y(n13763) );
  inv_1 U13190 ( .A(n13438), .Y(n13582) );
  nand2_1 U13191 ( .A(n13936), .B(n13910), .Y(n13438) );
  inv_1 U13192 ( .A(n13874), .Y(n13722) );
  inv_1 U13193 ( .A(n13937), .Y(n13752) );
  nand2_1 U13194 ( .A(n13920), .B(n13743), .Y(n13568) );
  nand2_1 U13195 ( .A(n13855), .B(n13920), .Y(n13488) );
  inv_1 U13196 ( .A(n13827), .Y(n13855) );
  inv_1 U13197 ( .A(n13853), .Y(n13553) );
  nor3_1 U13198 ( .A(n13827), .B(n13874), .C(n13825), .Y(n13853) );
  nand3_1 U13199 ( .A(n13886), .B(n12968), .C(n13938), .Y(n13825) );
  nand2_1 U13200 ( .A(n13931), .B(n13939), .Y(n13874) );
  nor2_1 U13201 ( .A(n13537), .B(n13524), .Y(n13902) );
  nand3_1 U13202 ( .A(n13846), .B(n13850), .C(n13786), .Y(n13524) );
  inv_1 U13203 ( .A(n13817), .Y(n13846) );
  nand3_1 U13204 ( .A(n13845), .B(n13940), .C(n23903), .Y(n13817) );
  nor4_1 U13205 ( .A(n13804), .B(n13663), .C(n13700), .D(n13797), .Y(n13878)
         );
  o221ai_1 U13206 ( .A1(n13475), .A2(n13476), .B1(n13483), .B2(n13635), .C1(
        n13941), .Y(n13797) );
  a21oi_1 U13207 ( .A1(n13717), .A2(n13510), .B1(n13942), .Y(n13941) );
  inv_1 U13208 ( .A(n13675), .Y(n13942) );
  nand2_1 U13209 ( .A(n13456), .B(n13439), .Y(n13675) );
  inv_1 U13210 ( .A(n13602), .Y(n13439) );
  nand2_1 U13211 ( .A(n13917), .B(n13936), .Y(n13602) );
  inv_1 U13212 ( .A(n13723), .Y(n13456) );
  nand3_1 U13213 ( .A(n13724), .B(n13721), .C(n13884), .Y(n13723) );
  nor2_1 U13214 ( .A(n13943), .B(n13944), .Y(n13724) );
  inv_1 U13215 ( .A(n13537), .Y(n13510) );
  nand2_1 U13216 ( .A(n13945), .B(n13911), .Y(n13537) );
  inv_1 U13217 ( .A(n12606), .Y(n13717) );
  nand2_1 U13218 ( .A(n13870), .B(n13843), .Y(n12606) );
  nor2_1 U13219 ( .A(n13946), .B(n23903), .Y(n13843) );
  and2_0 U13220 ( .A(n13835), .B(n13837), .X(n13870) );
  nor2_1 U13221 ( .A(n13947), .B(n13948), .Y(n13835) );
  inv_1 U13222 ( .A(n12568), .Y(n13635) );
  o21ai_0 U13223 ( .A1(n13945), .A2(n12599), .B1(n13918), .Y(n12568) );
  a21oi_1 U13224 ( .A1(n13625), .A2(n13626), .B1(n13509), .Y(n13483) );
  inv_1 U13225 ( .A(n12592), .Y(n13509) );
  nand2_1 U13226 ( .A(n13720), .B(n13920), .Y(n12592) );
  inv_1 U13227 ( .A(n13898), .Y(n13720) );
  inv_1 U13228 ( .A(n13873), .Y(n13626) );
  nand2_1 U13229 ( .A(n13820), .B(n13938), .Y(n13873) );
  nor2_1 U13230 ( .A(n13764), .B(n13827), .Y(n13625) );
  nand2_1 U13231 ( .A(n13915), .B(n13921), .Y(n13827) );
  nand2_1 U13232 ( .A(n13891), .B(n13892), .Y(n13476) );
  and2_0 U13233 ( .A(n13838), .B(n13833), .X(n13892) );
  and2_0 U13234 ( .A(n13935), .B(n13938), .X(n13891) );
  inv_1 U13235 ( .A(n13672), .Y(n13475) );
  o21ai_0 U13236 ( .A1(n13949), .A2(n12599), .B1(n13925), .Y(n13672) );
  o211ai_1 U13237 ( .A1(n12596), .A2(n12594), .B1(n13739), .C1(n13453), .Y(
        n13700) );
  nand2_1 U13238 ( .A(n13620), .B(n12569), .Y(n13453) );
  and3_1 U13239 ( .A(n13743), .B(n13830), .C(n13721), .X(n12569) );
  and2_0 U13240 ( .A(n13820), .B(n13885), .X(n13721) );
  nor2_1 U13241 ( .A(n13950), .B(n23903), .Y(n13820) );
  nor2_1 U13242 ( .A(n13943), .B(n13951), .Y(n13830) );
  nand4_1 U13243 ( .A(n13741), .B(n13742), .C(n13458), .D(n13725), .Y(n13739)
         );
  inv_1 U13244 ( .A(n13756), .Y(n13458) );
  inv_1 U13245 ( .A(n13828), .Y(n13742) );
  nand3_1 U13246 ( .A(n13924), .B(n12968), .C(n13938), .Y(n13828) );
  inv_1 U13247 ( .A(n13429), .Y(n12594) );
  nand2_1 U13248 ( .A(n12757), .B(n13736), .Y(n13429) );
  nand2_1 U13249 ( .A(n13893), .B(n13838), .Y(n13736) );
  and2_0 U13250 ( .A(n13895), .B(n13841), .X(n13893) );
  and3_1 U13251 ( .A(n23990), .B(n12968), .C(n13952), .X(n13841) );
  and2_0 U13252 ( .A(n13931), .B(n13845), .X(n13895) );
  inv_1 U13253 ( .A(n13460), .Y(n12596) );
  o21ai_0 U13254 ( .A1(n13945), .A2(n12599), .B1(n13925), .Y(n13460) );
  o221ai_1 U13255 ( .A1(n13472), .A2(n13575), .B1(n13756), .B2(n13789), .C1(
        n13953), .Y(n13663) );
  a21oi_1 U13256 ( .A1(n13788), .A2(n13442), .B1(n13623), .Y(n13953) );
  and3_1 U13257 ( .A(n13920), .B(n13620), .C(n13884), .X(n13623) );
  inv_1 U13258 ( .A(n12593), .Y(n13620) );
  nand2_1 U13259 ( .A(n13936), .B(n13945), .Y(n12593) );
  nor2_1 U13260 ( .A(n13954), .B(inData[27]), .Y(n13945) );
  and3_1 U13261 ( .A(n13935), .B(n13885), .C(n13848), .X(n13920) );
  inv_1 U13262 ( .A(n13955), .Y(n13848) );
  o21ai_0 U13263 ( .A1(n13949), .A2(n12599), .B1(n13918), .Y(n13442) );
  inv_1 U13264 ( .A(n13427), .Y(n13788) );
  nand2_1 U13265 ( .A(n13834), .B(n13783), .Y(n13427) );
  inv_1 U13266 ( .A(n13818), .Y(n13783) );
  nand4_1 U13267 ( .A(n13885), .B(n13867), .C(n13886), .D(n13868), .Y(n13818)
         );
  nand2_1 U13268 ( .A(n13909), .B(n13832), .Y(n13789) );
  and2_0 U13269 ( .A(n13860), .B(n13831), .X(n13909) );
  nand2_1 U13270 ( .A(n13949), .B(n13936), .Y(n13756) );
  inv_1 U13271 ( .A(n13925), .Y(n13936) );
  nand3_1 U13272 ( .A(n13786), .B(n13850), .C(n13834), .Y(n13575) );
  nor3_1 U13273 ( .A(n13956), .B(n13944), .C(n12968), .Y(n13834) );
  and2_0 U13274 ( .A(n13926), .B(n13868), .X(n13850) );
  nor3_1 U13275 ( .A(n13928), .B(n13929), .C(n13957), .Y(n13786) );
  inv_1 U13276 ( .A(n13512), .Y(n13472) );
  o21ai_0 U13277 ( .A1(n13910), .A2(n12599), .B1(n13925), .Y(n13512) );
  nand2_1 U13278 ( .A(n12574), .B(n13958), .Y(n13925) );
  inv_1 U13279 ( .A(n12574), .Y(n12599) );
  nor2_1 U13280 ( .A(n13959), .B(n13954), .Y(n13910) );
  o21ai_0 U13281 ( .A1(n13446), .A2(n13584), .B1(n13744), .Y(n13804) );
  or4_1 U13282 ( .A(n13858), .B(n13764), .C(n13960), .D(n13947), .X(n13744) );
  nand3_1 U13283 ( .A(n13935), .B(n13885), .C(n12615), .Y(n13858) );
  inv_1 U13284 ( .A(n13648), .Y(n12615) );
  nand2_1 U13285 ( .A(n13917), .B(n13911), .Y(n13648) );
  nor2_1 U13286 ( .A(inData[27]), .B(inData[31]), .Y(n13917) );
  nor2_1 U13287 ( .A(n13957), .B(n23903), .Y(n13935) );
  nand3_1 U13288 ( .A(n13836), .B(n13833), .C(n13859), .Y(n13584) );
  inv_1 U13289 ( .A(n13961), .Y(n13859) );
  nor2_1 U13290 ( .A(n13962), .B(n23903), .Y(n13836) );
  nand2_1 U13291 ( .A(n13949), .B(n13911), .Y(n13446) );
  inv_1 U13292 ( .A(n13918), .Y(n13911) );
  nand2_1 U13293 ( .A(inData[17]), .B(n12574), .Y(n13918) );
  nand3_1 U13294 ( .A(n13354), .B(n13351), .C(n13275), .Y(n12574) );
  and2_0 U13295 ( .A(n13387), .B(n13397), .X(n13354) );
  nor2_1 U13296 ( .A(n13959), .B(inData[31]), .Y(n13949) );
  o221ai_1 U13297 ( .A1(n13963), .A2(n12747), .B1(n13964), .B2(n10683), .C1(
        n13965), .Y(n10398) );
  o21ai_0 U13298 ( .A1(n13966), .A2(n13967), .B1(n10685), .Y(n13965) );
  nand4_1 U13299 ( .A(n13968), .B(n13969), .C(n13970), .D(n13971), .Y(n13967)
         );
  nor3_1 U13300 ( .A(n13972), .B(n10705), .C(n13973), .Y(n13971) );
  nand4_1 U13301 ( .A(n13974), .B(n13975), .C(n13976), .D(n13977), .Y(n13966)
         );
  and3_1 U13302 ( .A(n13978), .B(n13979), .C(n10719), .X(n13977) );
  nor4_1 U13303 ( .A(n13980), .B(n13981), .C(n13982), .D(n13983), .Y(n13964)
         );
  nand3_1 U13304 ( .A(n13984), .B(n13985), .C(n13986), .Y(n13981) );
  nand4_1 U13305 ( .A(n13987), .B(n10694), .C(n13988), .D(n13989), .Y(n13980)
         );
  nor2_1 U13306 ( .A(n13990), .B(n13991), .Y(n13989) );
  nor4_1 U13307 ( .A(n13992), .B(n13993), .C(n13994), .D(n13995), .Y(n13963)
         );
  nand3_1 U13308 ( .A(n10699), .B(n10695), .C(n13996), .Y(n13993) );
  or4_1 U13309 ( .A(n13997), .B(n13998), .C(n12781), .D(n12764), .X(n13992) );
  nand4_1 U13310 ( .A(n13999), .B(n14000), .C(n14001), .D(n14002), .Y(n12764)
         );
  and4_1 U13311 ( .A(n14003), .B(n14004), .C(n14005), .D(n14006), .X(n14002)
         );
  nand3_1 U13312 ( .A(n14007), .B(n10696), .C(n14008), .Y(n12781) );
  o211ai_1 U13313 ( .A1(n14009), .A2(n10683), .B1(n14010), .C1(n14011), .Y(
        n10397) );
  o21ai_0 U13314 ( .A1(n14012), .A2(n14013), .B1(n12757), .Y(n14011) );
  nand4_1 U13315 ( .A(n14014), .B(n14015), .C(n14016), .D(n14017), .Y(n14013)
         );
  inv_1 U13316 ( .A(n13998), .Y(n14014) );
  nand3_1 U13317 ( .A(n10701), .B(n10709), .C(n12777), .Y(n13998) );
  nand4_1 U13318 ( .A(n14001), .B(n14018), .C(n10725), .D(n14019), .Y(n14012)
         );
  o21ai_0 U13319 ( .A1(n14020), .A2(n14021), .B1(n10685), .Y(n14010) );
  nand4_1 U13320 ( .A(n14022), .B(n14023), .C(n12774), .D(n14006), .Y(n14021)
         );
  nand4_1 U13321 ( .A(n14024), .B(n10692), .C(n10693), .D(n14025), .Y(n14020)
         );
  nor4_1 U13322 ( .A(n14026), .B(n14027), .C(n14028), .D(n13994), .Y(n14009)
         );
  nand3_1 U13323 ( .A(n10718), .B(n13979), .C(n14029), .Y(n14027) );
  nand4_1 U13324 ( .A(n14030), .B(n14031), .C(n14032), .D(n14033), .Y(n14026)
         );
  o211ai_1 U13325 ( .A1(n14034), .A2(n10683), .B1(n14035), .C1(n14036), .Y(
        n10396) );
  o21ai_0 U13326 ( .A1(n14037), .A2(n14038), .B1(n10685), .Y(n14036) );
  nand4_1 U13327 ( .A(n14039), .B(n14022), .C(n13984), .D(n14040), .Y(n14038)
         );
  inv_1 U13328 ( .A(n14041), .Y(n13984) );
  nor3_1 U13329 ( .A(n14042), .B(n14043), .C(n14044), .Y(n14022) );
  inv_1 U13330 ( .A(n14045), .Y(n14043) );
  nand4_1 U13331 ( .A(n14000), .B(n14003), .C(n14046), .D(n10701), .Y(n14037)
         );
  o21ai_0 U13332 ( .A1(n14047), .A2(n14048), .B1(n12757), .Y(n14035) );
  nand4_1 U13333 ( .A(n14049), .B(n14032), .C(n14017), .D(n14050), .Y(n14048)
         );
  and3_1 U13334 ( .A(n14051), .B(n10720), .C(n14052), .X(n14032) );
  nand4_1 U13335 ( .A(n10719), .B(n14024), .C(n12777), .D(n10695), .Y(n14047)
         );
  nor4_1 U13336 ( .A(n14053), .B(n14054), .C(n12765), .D(n14055), .Y(n14034)
         );
  nand3_1 U13337 ( .A(n14056), .B(n14057), .C(n10725), .Y(n14054) );
  nand4_1 U13338 ( .A(n14058), .B(n14059), .C(n14030), .D(n14060), .Y(n14053)
         );
  and4_1 U13339 ( .A(n14061), .B(n14062), .C(n14063), .D(n14064), .X(n14030)
         );
  and4_1 U13340 ( .A(n14065), .B(n13975), .C(n12772), .D(n14066), .X(n14064)
         );
  inv_1 U13341 ( .A(n12769), .Y(n14066) );
  nor2_1 U13342 ( .A(n14067), .B(n14068), .Y(n14063) );
  inv_1 U13343 ( .A(n14069), .Y(n14059) );
  o211ai_1 U13344 ( .A1(n14070), .A2(n10683), .B1(n14071), .C1(n14072), .Y(
        n10395) );
  o21ai_0 U13345 ( .A1(n14073), .A2(n14074), .B1(n12757), .Y(n14072) );
  or4_1 U13346 ( .A(n14075), .B(n14076), .C(n13973), .D(n13997), .X(n14074) );
  nand3_1 U13347 ( .A(n14077), .B(n14024), .C(n14078), .Y(n13973) );
  nand4_1 U13348 ( .A(n14079), .B(n14001), .C(n14080), .D(n14081), .Y(n14073)
         );
  inv_1 U13349 ( .A(n14082), .Y(n14079) );
  o21ai_0 U13350 ( .A1(n14083), .A2(n14084), .B1(n10685), .Y(n14071) );
  nand4_1 U13351 ( .A(n14085), .B(n14086), .C(n14087), .D(n14088), .Y(n14084)
         );
  nor3_1 U13352 ( .A(n12785), .B(n14055), .C(n10691), .Y(n14088) );
  inv_1 U13353 ( .A(n14089), .Y(n14087) );
  nand4_1 U13354 ( .A(n14004), .B(n14090), .C(n14000), .D(n14091), .Y(n14083)
         );
  and3_1 U13355 ( .A(n14092), .B(n12777), .C(n14093), .X(n14091) );
  nor4_1 U13356 ( .A(n14094), .B(n14095), .C(n10722), .D(n14096), .Y(n14070)
         );
  nand3_1 U13357 ( .A(n14097), .B(n14061), .C(n14098), .Y(n14095) );
  or4_1 U13358 ( .A(n14099), .B(n14100), .C(n13983), .D(n12769), .X(n14094) );
  nand4_1 U13359 ( .A(n14101), .B(n10727), .C(n14102), .D(n14103), .Y(n12769)
         );
  and2_0 U13360 ( .A(n13974), .B(n13976), .X(n14103) );
  nand4_1 U13361 ( .A(n14104), .B(n10718), .C(n14060), .D(n14105), .Y(n13983)
         );
  nor4_1 U13362 ( .A(n14106), .B(n12844), .C(n14107), .D(n10716), .Y(n14105)
         );
  inv_1 U13363 ( .A(n14108), .Y(n10716) );
  o221ai_1 U13364 ( .A1(n14109), .A2(n10683), .B1(n14110), .B2(n12750), .C1(
        n14111), .Y(n10394) );
  o21ai_0 U13365 ( .A1(n14112), .A2(n14113), .B1(n12757), .Y(n14111) );
  nand4_1 U13366 ( .A(n14114), .B(n14115), .C(n14116), .D(n14016), .Y(n14113)
         );
  nand4_1 U13367 ( .A(n14117), .B(n14078), .C(n10706), .D(n12777), .Y(n14112)
         );
  nor4_1 U13368 ( .A(n14118), .B(n14119), .C(n14120), .D(n14121), .Y(n14110)
         );
  nand3_1 U13369 ( .A(n14023), .B(n12774), .C(n14122), .Y(n14119) );
  inv_1 U13370 ( .A(n10723), .Y(n14023) );
  nand3_1 U13371 ( .A(n14123), .B(n12751), .C(n14124), .Y(n14118) );
  and3_1 U13372 ( .A(n10725), .B(n12778), .C(n14019), .X(n14124) );
  nor4_1 U13373 ( .A(n14125), .B(n14126), .C(n14127), .D(n14068), .Y(n14109)
         );
  inv_1 U13374 ( .A(n14004), .Y(n14068) );
  inv_1 U13375 ( .A(n14101), .Y(n14127) );
  nand3_1 U13376 ( .A(n14062), .B(n10693), .C(n14108), .Y(n14126) );
  or4_1 U13377 ( .A(n14128), .B(n14129), .C(n14130), .D(n13991), .X(n14125) );
  o21ai_0 U13378 ( .A1(n14131), .A2(n12747), .B1(n14132), .Y(n10393) );
  mux2i_1 U13379 ( .A0(n10685), .A1(n14133), .S(n14134), .Y(n14132) );
  nor4_1 U13380 ( .A(n14135), .B(n14136), .C(n14041), .D(n14100), .Y(n14134)
         );
  nand2_1 U13381 ( .A(n14137), .B(n14138), .Y(n14041) );
  nand4_1 U13382 ( .A(n14114), .B(n14139), .C(n14033), .D(n13979), .Y(n14135)
         );
  nor4_1 U13383 ( .A(n14140), .B(n14141), .C(n10683), .D(n14142), .Y(n14133)
         );
  nand2_1 U13384 ( .A(n14016), .B(n14143), .Y(n14142) );
  nand3_1 U13385 ( .A(n14144), .B(n14031), .C(n14145), .Y(n14141) );
  and4_1 U13386 ( .A(n14108), .B(n10708), .C(n14117), .D(n14146), .X(n14031)
         );
  nor2_1 U13387 ( .A(n13991), .B(n14147), .Y(n14146) );
  inv_1 U13388 ( .A(n14148), .Y(n14144) );
  nand4_1 U13389 ( .A(n14102), .B(n14005), .C(n13974), .D(n14149), .Y(n14140)
         );
  and4_1 U13390 ( .A(n14024), .B(n10717), .C(n14056), .D(n14101), .X(n14149)
         );
  nor4_1 U13391 ( .A(n14150), .B(n14151), .C(n12766), .D(n14152), .Y(n14131)
         );
  inv_1 U13392 ( .A(n13987), .Y(n14152) );
  nand3_1 U13393 ( .A(n14153), .B(n10710), .C(n14081), .Y(n14151) );
  nand3_1 U13394 ( .A(n14154), .B(n14122), .C(n14155), .Y(n14150) );
  nor3_1 U13395 ( .A(n14128), .B(n14156), .C(n12765), .Y(n14155) );
  inv_1 U13396 ( .A(n13988), .Y(n12765) );
  nand4_1 U13397 ( .A(n13976), .B(n14157), .C(n14006), .D(n13978), .Y(n14128)
         );
  and3_1 U13398 ( .A(n13975), .B(n10718), .C(n13985), .X(n14122) );
  inv_1 U13399 ( .A(n14158), .Y(n14154) );
  o221ai_1 U13400 ( .A1(n14159), .A2(n12747), .B1(n14160), .B2(n12750), .C1(
        n14161), .Y(n10392) );
  o21ai_0 U13401 ( .A1(n14162), .A2(n14163), .B1(n14164), .Y(n14161) );
  or4_1 U13402 ( .A(n14120), .B(n14129), .C(n10724), .D(n14165), .X(n14163) );
  nand4_1 U13403 ( .A(n14166), .B(n14101), .C(n14167), .D(n14168), .Y(n10724)
         );
  nor4_1 U13404 ( .A(n12766), .B(n14067), .C(n14169), .D(n14170), .Y(n14168)
         );
  inv_1 U13405 ( .A(n13978), .Y(n14067) );
  inv_1 U13406 ( .A(n14097), .Y(n12766) );
  and3_1 U13407 ( .A(n12751), .B(n14171), .C(n14081), .X(n14167) );
  nand3_1 U13408 ( .A(n10701), .B(n10708), .C(n14172), .Y(n14129) );
  nand4_1 U13409 ( .A(n14017), .B(n14045), .C(n14173), .D(n10720), .Y(n14120)
         );
  and2_0 U13410 ( .A(n10709), .B(n13979), .X(n14173) );
  nand4_1 U13411 ( .A(n10710), .B(n14025), .C(n10707), .D(n14174), .Y(n14162)
         );
  and2_0 U13412 ( .A(n14024), .B(n14060), .X(n14174) );
  nor4_1 U13413 ( .A(n14175), .B(n14176), .C(n14042), .D(n14076), .Y(n14160)
         );
  nand3_1 U13414 ( .A(n14177), .B(n14178), .C(n13985), .Y(n14042) );
  nand3_1 U13415 ( .A(n13969), .B(n13976), .C(n14179), .Y(n14176) );
  nand4_1 U13416 ( .A(n14180), .B(n10693), .C(n14123), .D(n14181), .Y(n14175)
         );
  and3_1 U13417 ( .A(n14033), .B(n13988), .C(n14117), .X(n14181) );
  nor4_1 U13418 ( .A(n14182), .B(n14183), .C(n14158), .D(n14136), .Y(n14159)
         );
  nand3_1 U13419 ( .A(n14029), .B(n14004), .C(n12772), .Y(n14136) );
  nand4_1 U13420 ( .A(n14001), .B(n14078), .C(n14184), .D(n14185), .Y(n14158)
         );
  and3_1 U13421 ( .A(n14186), .B(n14092), .C(n14003), .X(n14185) );
  and3_1 U13422 ( .A(n10692), .B(n10699), .C(n14062), .X(n14186) );
  and3_1 U13423 ( .A(n14051), .B(n14187), .C(n14065), .X(n14184) );
  nand3_1 U13424 ( .A(n14015), .B(n14188), .C(n14189), .Y(n14183) );
  nand4_1 U13425 ( .A(n14040), .B(n14007), .C(n14190), .D(n14080), .Y(n14182)
         );
  and2_0 U13426 ( .A(n10700), .B(n14093), .X(n14190) );
  o221ai_1 U13427 ( .A1(n14191), .A2(n12747), .B1(n14192), .B2(n10683), .C1(
        n14193), .Y(n10391) );
  o21ai_0 U13428 ( .A1(n14194), .A2(n14195), .B1(n10685), .Y(n14193) );
  nand4_1 U13429 ( .A(n14145), .B(n14058), .C(n14008), .D(n14138), .Y(n14195)
         );
  inv_1 U13430 ( .A(n14096), .Y(n14008) );
  nand2_1 U13431 ( .A(n14029), .B(n10726), .Y(n14096) );
  nor3_1 U13432 ( .A(n14196), .B(n12844), .C(n14075), .Y(n14058) );
  nand4_1 U13433 ( .A(n13979), .B(n10696), .C(n14006), .D(n14197), .Y(n14075)
         );
  and3_1 U13434 ( .A(n14117), .B(n14007), .C(n13999), .X(n14197) );
  and3_1 U13435 ( .A(n14017), .B(n14057), .C(n13970), .X(n14145) );
  nand4_1 U13436 ( .A(n14097), .B(n10694), .C(n12775), .D(n14046), .Y(n14194)
         );
  nor4_1 U13437 ( .A(n14198), .B(n14199), .C(n14200), .D(n14156), .Y(n14192)
         );
  inv_1 U13438 ( .A(n14171), .Y(n14200) );
  nand3_1 U13439 ( .A(n10695), .B(n10708), .C(n10717), .Y(n14199) );
  or4_1 U13440 ( .A(n14099), .B(n13982), .C(n13997), .D(n14201), .X(n14198) );
  nand3_1 U13441 ( .A(n10710), .B(n14025), .C(n14123), .Y(n13997) );
  nand3_1 U13442 ( .A(n12773), .B(n14081), .C(n14189), .Y(n13982) );
  and3_1 U13443 ( .A(n14050), .B(n12774), .C(n12759), .X(n14189) );
  nand3_1 U13444 ( .A(n10720), .B(n10719), .C(n14018), .Y(n14099) );
  nor4_1 U13445 ( .A(n14202), .B(n14203), .C(n12763), .D(n14100), .Y(n14191)
         );
  nand2_1 U13446 ( .A(n10701), .B(n12778), .Y(n14100) );
  nand3_1 U13447 ( .A(n14204), .B(n14137), .C(n14205), .Y(n14203) );
  nand4_1 U13448 ( .A(n14005), .B(n14056), .C(n14206), .D(n14077), .Y(n14202)
         );
  and2_0 U13449 ( .A(n14207), .B(n14153), .X(n14206) );
  o221ai_1 U13450 ( .A1(n14208), .A2(n10683), .B1(n12747), .B2(n14209), .C1(
        n14210), .Y(n10390) );
  o21ai_0 U13451 ( .A1(n14211), .A2(n14212), .B1(n10685), .Y(n14210) );
  nand4_1 U13452 ( .A(n14213), .B(n14214), .C(n14049), .D(n14086), .Y(n14212)
         );
  inv_1 U13453 ( .A(n14044), .Y(n14086) );
  o21ai_0 U13454 ( .A1(n14215), .A2(n14216), .B1(n12759), .Y(n14044) );
  and4_1 U13455 ( .A(n14217), .B(n14218), .C(n14093), .D(n10692), .X(n14049)
         );
  inv_1 U13456 ( .A(n14076), .Y(n14217) );
  nand3_1 U13457 ( .A(n12760), .B(n14219), .C(n14116), .Y(n14076) );
  inv_1 U13458 ( .A(n14220), .Y(n14214) );
  nand4_1 U13459 ( .A(n14157), .B(n14123), .C(n14221), .D(n10710), .Y(n14211)
         );
  nor3_1 U13460 ( .A(n14222), .B(n12752), .C(n14223), .Y(n14209) );
  nand3_1 U13461 ( .A(n14138), .B(n14005), .C(n14204), .Y(n14222) );
  nor4_1 U13462 ( .A(n14224), .B(n14121), .C(n14225), .D(n14170), .Y(n14208)
         );
  nand4_1 U13463 ( .A(n14153), .B(n10700), .C(n14024), .D(n14226), .Y(n14121)
         );
  nor3_1 U13464 ( .A(n13995), .B(n14107), .C(n13994), .Y(n14226) );
  inv_1 U13465 ( .A(n14080), .Y(n13994) );
  inv_1 U13466 ( .A(n12775), .Y(n14107) );
  nand3_1 U13467 ( .A(n14187), .B(n12777), .C(n14227), .Y(n14224) );
  o21ai_0 U13468 ( .A1(n14228), .A2(n10683), .B1(n14229), .Y(n10389) );
  mux2i_1 U13469 ( .A0(n10685), .A1(n14230), .S(n14231), .Y(n14229) );
  nor4_1 U13470 ( .A(n14232), .B(n14233), .C(n14089), .D(n14148), .Y(n14231)
         );
  nand3_1 U13471 ( .A(n14052), .B(n13988), .C(n14234), .Y(n14089) );
  inv_1 U13472 ( .A(n12770), .Y(n14234) );
  nand3_1 U13473 ( .A(n14062), .B(n10699), .C(n14017), .Y(n12770) );
  nand3_1 U13474 ( .A(n14235), .B(n13999), .C(n14236), .Y(n14233) );
  inv_1 U13475 ( .A(n13972), .Y(n14236) );
  nand4_1 U13476 ( .A(n14033), .B(n14065), .C(n14221), .D(n14180), .Y(n13972)
         );
  nand4_1 U13477 ( .A(n10694), .B(n10697), .C(n10725), .D(n14237), .Y(n14232)
         );
  and3_1 U13478 ( .A(n14018), .B(n14051), .C(n14098), .X(n14237) );
  nor4_1 U13479 ( .A(n14238), .B(n14239), .C(n10704), .D(n14240), .Y(n14230)
         );
  nand3_1 U13480 ( .A(n14143), .B(n14005), .C(n14241), .Y(n10704) );
  and3_1 U13481 ( .A(n14004), .B(n12757), .C(n14104), .X(n14241) );
  nand3_1 U13482 ( .A(n12783), .B(n14204), .C(n14015), .Y(n14239) );
  inv_1 U13483 ( .A(n14242), .Y(n14015) );
  inv_1 U13484 ( .A(n12752), .Y(n12783) );
  nand4_1 U13485 ( .A(n14123), .B(n14101), .C(n14006), .D(n14243), .Y(n14238)
         );
  nor2_1 U13486 ( .A(n14156), .B(n14244), .Y(n14243) );
  inv_1 U13487 ( .A(n14000), .Y(n14156) );
  inv_1 U13488 ( .A(n14240), .Y(n14228) );
  nand4_1 U13489 ( .A(n14218), .B(n14245), .C(n14246), .D(n14247), .Y(n14240)
         );
  and4_1 U13490 ( .A(n10719), .B(n10727), .C(n14166), .D(n13978), .X(n14247)
         );
  nor2_1 U13491 ( .A(n14248), .B(n14249), .Y(n14246) );
  inv_1 U13492 ( .A(n13986), .Y(n14249) );
  nor3_1 U13493 ( .A(n14250), .B(n14196), .C(n14170), .Y(n13986) );
  inv_1 U13494 ( .A(n10700), .Y(n14196) );
  inv_1 U13495 ( .A(n14092), .Y(n14250) );
  o221ai_1 U13496 ( .A1(n14251), .A2(n12750), .B1(n14252), .B2(n10683), .C1(
        n14253), .Y(n10388) );
  o21ai_0 U13497 ( .A1(n14254), .A2(n14255), .B1(n12757), .Y(n14253) );
  nand4_1 U13498 ( .A(n14213), .B(n14256), .C(n13970), .D(n12772), .Y(n14255)
         );
  inv_1 U13499 ( .A(n10722), .Y(n13970) );
  inv_1 U13500 ( .A(n12780), .Y(n14256) );
  nand4_1 U13501 ( .A(n14033), .B(n14178), .C(n14138), .D(n14257), .Y(n12780)
         );
  and4_1 U13502 ( .A(n14093), .B(n14092), .C(n10720), .D(n14018), .X(n14257)
         );
  and4_1 U13503 ( .A(n14004), .B(n14003), .C(n14062), .D(n13979), .X(n14213)
         );
  nand4_1 U13504 ( .A(n13974), .B(n12760), .C(n14001), .D(n14153), .Y(n14254)
         );
  nor4_1 U13505 ( .A(n14258), .B(n14259), .C(n14260), .D(n14261), .Y(n14252)
         );
  nand4_1 U13506 ( .A(n14039), .B(n14235), .C(n13985), .D(n14102), .Y(n14261)
         );
  inv_1 U13507 ( .A(n12763), .Y(n14235) );
  nand3_1 U13508 ( .A(n14080), .B(n10718), .C(n14172), .Y(n12763) );
  nor3_1 U13509 ( .A(n14028), .B(n14262), .C(n14242), .Y(n14039) );
  inv_1 U13510 ( .A(n14123), .Y(n14028) );
  nand4_1 U13511 ( .A(n13975), .B(n13988), .C(n14104), .D(n14187), .Y(n14260)
         );
  nand4_1 U13512 ( .A(n12751), .B(n10694), .C(n14024), .D(n12777), .Y(n14259)
         );
  nand4_1 U13513 ( .A(n10692), .B(n14057), .C(n10707), .D(n14263), .Y(n14258)
         );
  nor4_1 U13514 ( .A(n14264), .B(n14265), .C(n14220), .D(n14266), .Y(n14251)
         );
  nand3_1 U13515 ( .A(n10709), .B(n14267), .C(n14040), .Y(n14220) );
  nand3_1 U13516 ( .A(n14268), .B(n14006), .C(n14085), .Y(n14265) );
  and3_1 U13517 ( .A(n14056), .B(n10693), .C(n13978), .X(n14085) );
  inv_1 U13518 ( .A(n12782), .Y(n14268) );
  nand4_1 U13519 ( .A(n14050), .B(n14177), .C(n14052), .D(n14269), .Y(n12782)
         );
  nor3_1 U13520 ( .A(n13991), .B(n14270), .C(n13990), .Y(n14269) );
  inv_1 U13521 ( .A(n14219), .Y(n13991) );
  nand4_1 U13522 ( .A(n14077), .B(n12778), .C(n10725), .D(n14271), .Y(n14264)
         );
  and2_0 U13523 ( .A(n14065), .B(n14051), .X(n14271) );
  o211ai_1 U13524 ( .A1(n14272), .A2(n12844), .B1(n14273), .C1(n14274), .Y(
        n10387) );
  o21ai_0 U13525 ( .A1(n14275), .A2(n14276), .B1(n10749), .Y(n14274) );
  nand4_1 U13526 ( .A(n14277), .B(n14278), .C(n14279), .D(n14280), .Y(n14276)
         );
  nor3_1 U13527 ( .A(n14281), .B(n14282), .C(n14283), .Y(n14280) );
  nand4_1 U13528 ( .A(n14284), .B(n14285), .C(n14286), .D(n14287), .Y(n14275)
         );
  nor4_1 U13529 ( .A(n14288), .B(n14289), .C(n14290), .D(n10767), .Y(n14287)
         );
  o21ai_0 U13530 ( .A1(n14291), .A2(n14292), .B1(n12847), .Y(n14273) );
  nand4_1 U13531 ( .A(n14293), .B(n14294), .C(n14295), .D(n14296), .Y(n14292)
         );
  a211oi_1 U13532 ( .A1(n14297), .A2(n14298), .B1(n12851), .C1(n14299), .Y(
        n14296) );
  inv_1 U13533 ( .A(n14300), .Y(n14295) );
  nand4_1 U13534 ( .A(n14301), .B(n14302), .C(n14303), .D(n14304), .Y(n14291)
         );
  and4_1 U13535 ( .A(n14305), .B(n14306), .C(n14307), .D(n14308), .X(n14304)
         );
  nor4_1 U13536 ( .A(n14309), .B(n14310), .C(n14311), .D(n14312), .Y(n14272)
         );
  nand3_1 U13537 ( .A(n14313), .B(n14314), .C(n14315), .Y(n14310) );
  nand4_1 U13538 ( .A(n14316), .B(n14317), .C(n14318), .D(n14319), .Y(n14309)
         );
  and2_0 U13539 ( .A(n14320), .B(n14321), .X(n14318) );
  o221ai_1 U13540 ( .A1(n14322), .A2(n12842), .B1(n14323), .B2(n10747), .C1(
        n14324), .Y(n10386) );
  o21ai_0 U13541 ( .A1(n14325), .A2(n14326), .B1(n10697), .Y(n14324) );
  nand4_1 U13542 ( .A(n14327), .B(n14328), .C(n14329), .D(n14330), .Y(n14326)
         );
  and3_1 U13543 ( .A(n14331), .B(n14332), .C(n14316), .X(n14330) );
  nand4_1 U13544 ( .A(n14333), .B(n14305), .C(n14334), .D(n14335), .Y(n14325)
         );
  and3_1 U13545 ( .A(n14284), .B(n14336), .C(n14308), .X(n14335) );
  nor4_1 U13546 ( .A(n14337), .B(n14338), .C(n14339), .D(n14340), .Y(n14323)
         );
  nand3_1 U13547 ( .A(n14341), .B(n14342), .C(n14343), .Y(n14340) );
  nand4_1 U13548 ( .A(n14344), .B(n14345), .C(n14346), .D(n14347), .Y(n14339)
         );
  o211ai_1 U13549 ( .A1(n14348), .A2(n14349), .B1(n14350), .C1(n14351), .Y(
        n14338) );
  nand4_1 U13550 ( .A(n14352), .B(n14303), .C(n14353), .D(n14354), .Y(n14337)
         );
  nor4_1 U13551 ( .A(n14355), .B(n14356), .C(n14357), .D(n14311), .Y(n14322)
         );
  nand3_1 U13552 ( .A(n14358), .B(n14359), .C(n14360), .Y(n14311) );
  o211ai_1 U13553 ( .A1(n14361), .A2(n12848), .B1(n14362), .C1(n10759), .Y(
        n14356) );
  nand4_1 U13554 ( .A(n14301), .B(n14363), .C(n14364), .D(n14365), .Y(n14355)
         );
  and3_1 U13555 ( .A(n14366), .B(n14367), .C(n14368), .X(n14365) );
  o221ai_1 U13556 ( .A1(n14369), .A2(n12844), .B1(n14370), .B2(n10747), .C1(
        n14371), .Y(n10385) );
  o21ai_0 U13557 ( .A1(n14372), .A2(n14373), .B1(n10749), .Y(n14371) );
  nand4_1 U13558 ( .A(n14374), .B(n14343), .C(n14329), .D(n14375), .Y(n14373)
         );
  inv_1 U13559 ( .A(n14376), .Y(n14343) );
  inv_1 U13560 ( .A(n14377), .Y(n14374) );
  nand4_1 U13561 ( .A(n10761), .B(n10760), .C(n14378), .D(n14305), .Y(n14372)
         );
  nor4_1 U13562 ( .A(n14379), .B(n14380), .C(n14381), .D(n14382), .Y(n10760)
         );
  o21ai_0 U13563 ( .A1(n10757), .A2(n14348), .B1(n14362), .Y(n14382) );
  nor4_1 U13564 ( .A(n14383), .B(n14384), .C(n14385), .D(n14386), .Y(n14370)
         );
  nand4_1 U13565 ( .A(n14387), .B(n14353), .C(n14388), .D(n14389), .Y(n14383)
         );
  nor4_1 U13566 ( .A(n14390), .B(n14391), .C(n14392), .D(n14393), .Y(n14369)
         );
  inv_1 U13567 ( .A(n14394), .Y(n14393) );
  nand3_1 U13568 ( .A(n14333), .B(n14395), .C(n14302), .Y(n14391) );
  or4_1 U13569 ( .A(n14396), .B(n14397), .C(n14398), .D(n14282), .X(n14390) );
  o211ai_1 U13570 ( .A1(n14399), .A2(n12844), .B1(n14400), .C1(n14401), .Y(
        n10384) );
  mux2i_1 U13571 ( .A0(n10749), .A1(n14402), .S(n14403), .Y(n14401) );
  nor4_1 U13572 ( .A(n14404), .B(n14405), .C(n14281), .D(n14406), .Y(n14403)
         );
  nand3_1 U13573 ( .A(n14407), .B(n14408), .C(n14375), .Y(n14405) );
  inv_1 U13574 ( .A(n14409), .Y(n14407) );
  nand4_1 U13575 ( .A(n14305), .B(n14359), .C(n14354), .D(n14410), .Y(n14404)
         );
  and3_1 U13576 ( .A(n14316), .B(n14411), .C(n14351), .X(n14410) );
  nor4_1 U13577 ( .A(n14412), .B(n14413), .C(n14414), .D(n10747), .Y(n14402)
         );
  nand3_1 U13578 ( .A(n10766), .B(n14415), .C(n14331), .Y(n14413) );
  nand4_1 U13579 ( .A(n14333), .B(n14416), .C(n10757), .D(n14417), .Y(n14412)
         );
  nor2_1 U13580 ( .A(n14418), .B(n14419), .Y(n14417) );
  nor4_1 U13581 ( .A(n14420), .B(n14421), .C(n14357), .D(n14397), .Y(n14399)
         );
  nand3_1 U13582 ( .A(n14308), .B(n14422), .C(n14321), .Y(n14397) );
  nand3_1 U13583 ( .A(n14423), .B(n14424), .C(n14425), .Y(n14421) );
  nand4_1 U13584 ( .A(n10773), .B(n14334), .C(n10771), .D(n14426), .Y(n14420)
         );
  nor2_1 U13585 ( .A(n14379), .B(n14381), .Y(n14426) );
  o221ai_1 U13586 ( .A1(n14427), .A2(n12842), .B1(n14428), .B2(n10747), .C1(
        n14429), .Y(n10383) );
  o21ai_0 U13587 ( .A1(n14430), .A2(n14431), .B1(n10697), .Y(n14429) );
  nand4_1 U13588 ( .A(n14432), .B(n14329), .C(n14433), .D(n14434), .Y(n14431)
         );
  and4_1 U13589 ( .A(n14394), .B(n14423), .C(n14408), .D(n14435), .X(n14434)
         );
  inv_1 U13590 ( .A(n14436), .Y(n14433) );
  inv_1 U13591 ( .A(n14437), .Y(n14432) );
  nand4_1 U13592 ( .A(n14301), .B(n14358), .C(n14438), .D(n14439), .Y(n14430)
         );
  and4_1 U13593 ( .A(n14440), .B(n14333), .C(n14441), .D(n14321), .X(n14439)
         );
  nor4_1 U13594 ( .A(n14442), .B(n14443), .C(n14444), .D(n14283), .Y(n14428)
         );
  nand3_1 U13595 ( .A(n14445), .B(n14350), .C(n14314), .Y(n14443) );
  nand3_1 U13596 ( .A(n14446), .B(n14447), .C(n14448), .Y(n14442) );
  nor3_1 U13597 ( .A(n14449), .B(n14450), .C(n14379), .Y(n14448) );
  nor4_1 U13598 ( .A(n14451), .B(n14452), .C(n14453), .D(n14454), .Y(n14427)
         );
  a21oi_1 U13599 ( .A1(n14348), .A2(n10756), .B1(n10757), .Y(n14452) );
  o211ai_1 U13600 ( .A1(n14455), .A2(n14361), .B1(n14456), .C1(n14457), .Y(
        n14451) );
  o221ai_1 U13601 ( .A1(n14458), .A2(n12842), .B1(n14459), .B2(n10747), .C1(
        n14460), .Y(n10382) );
  o21ai_0 U13602 ( .A1(n14461), .A2(n14462), .B1(n10697), .Y(n14460) );
  or4_1 U13603 ( .A(n14312), .B(n14444), .C(n14463), .D(n14464), .X(n14462) );
  nand3_1 U13604 ( .A(n14351), .B(n14438), .C(n14352), .Y(n14464) );
  nand4_1 U13605 ( .A(n14345), .B(n14350), .C(n10772), .D(n14378), .Y(n14312)
         );
  nand4_1 U13606 ( .A(n14333), .B(n14354), .C(n14465), .D(n14466), .Y(n14461)
         );
  and3_1 U13607 ( .A(n14319), .B(n14308), .C(n14467), .X(n14466) );
  nor4_1 U13608 ( .A(n14468), .B(n14469), .C(n14357), .D(n14376), .Y(n14459)
         );
  nand3_1 U13609 ( .A(n14441), .B(n14470), .C(n14471), .Y(n14376) );
  o211ai_1 U13610 ( .A1(n14472), .A2(n14473), .B1(n14474), .C1(n14375), .Y(
        n14469) );
  nand4_1 U13611 ( .A(n14475), .B(n14306), .C(n14334), .D(n14476), .Y(n14468)
         );
  nor3_1 U13612 ( .A(n14419), .B(n14477), .C(n14290), .Y(n14476) );
  inv_1 U13613 ( .A(n14317), .Y(n14419) );
  nor2_1 U13614 ( .A(n14478), .B(n14479), .Y(n14458) );
  nand4_1 U13615 ( .A(n14480), .B(n14342), .C(n14481), .D(n14482), .Y(n14479)
         );
  and4_1 U13616 ( .A(n14286), .B(n14483), .C(n14423), .D(n14408), .X(n14482)
         );
  inv_1 U13617 ( .A(n14385), .Y(n14408) );
  and4_1 U13618 ( .A(n14424), .B(n14484), .C(n14320), .D(n14307), .X(n14342)
         );
  inv_1 U13619 ( .A(n14485), .Y(n14480) );
  nand4_1 U13620 ( .A(n14321), .B(n14302), .C(n14486), .D(n14487), .Y(n14478)
         );
  nor4_1 U13621 ( .A(n14488), .B(n14489), .C(n14490), .D(n14491), .Y(n14487)
         );
  inv_1 U13622 ( .A(n14416), .Y(n14488) );
  nand3_1 U13623 ( .A(n14492), .B(n14400), .C(n14493), .Y(n10381) );
  a22oi_1 U13624 ( .A1(n14494), .A2(n10697), .B1(n12847), .B2(n14495), .Y(
        n14493) );
  nand4_1 U13625 ( .A(n14303), .B(n14465), .C(n14496), .D(n14497), .Y(n14495)
         );
  and4_1 U13626 ( .A(n14424), .B(n14360), .C(n14341), .D(n14457), .X(n14497)
         );
  and3_1 U13627 ( .A(n14336), .B(n14498), .C(n14467), .X(n14457) );
  inv_1 U13628 ( .A(n14499), .Y(n14341) );
  nor3_1 U13629 ( .A(n14500), .B(n14288), .C(n14501), .Y(n14496) );
  inv_1 U13630 ( .A(n14378), .Y(n14500) );
  nand3_1 U13631 ( .A(n12843), .B(n14346), .C(n14502), .Y(n14494) );
  and3_1 U13632 ( .A(n14279), .B(n10765), .C(n14364), .X(n14502) );
  nor2_1 U13633 ( .A(n14503), .B(n14504), .Y(n12843) );
  inv_1 U13634 ( .A(n14358), .Y(n14504) );
  o21ai_0 U13635 ( .A1(n14505), .A2(n14506), .B1(n10749), .Y(n14492) );
  nand4_1 U13636 ( .A(n14507), .B(n14351), .C(n14314), .D(n14508), .Y(n14506)
         );
  nor3_1 U13637 ( .A(n14509), .B(n10764), .C(n14377), .Y(n14508) );
  nand3_1 U13638 ( .A(n14445), .B(n14316), .C(n10759), .Y(n14377) );
  nand4_1 U13639 ( .A(n14510), .B(n14306), .C(n14422), .D(n14511), .Y(n14505)
         );
  nor3_1 U13640 ( .A(n14512), .B(n10768), .C(n14290), .Y(n14511) );
  inv_1 U13641 ( .A(n14513), .Y(n14290) );
  o211ai_1 U13642 ( .A1(n12844), .A2(n14514), .B1(n14515), .C1(n14516), .Y(
        n10380) );
  o21ai_0 U13643 ( .A1(n14517), .A2(n14518), .B1(n12847), .Y(n14516) );
  or4_1 U13644 ( .A(n14384), .B(n14283), .C(n14509), .D(n14519), .X(n14518) );
  nand4_1 U13645 ( .A(n14285), .B(n14284), .C(n14352), .D(n14362), .Y(n14519)
         );
  nand3_1 U13646 ( .A(n14308), .B(n14363), .C(n14520), .Y(n14509) );
  and3_1 U13647 ( .A(n10771), .B(n14521), .C(n10772), .X(n14520) );
  nand4_1 U13648 ( .A(n14303), .B(n14366), .C(n14522), .D(n14354), .Y(n14384)
         );
  nor2_1 U13649 ( .A(n14523), .B(n14501), .Y(n14522) );
  nand4_1 U13650 ( .A(n14438), .B(n14524), .C(n14415), .D(n14525), .Y(n14517)
         );
  and4_1 U13651 ( .A(n14475), .B(n14334), .C(n14378), .D(n14358), .X(n14525)
         );
  inv_1 U13652 ( .A(n14526), .Y(n14475) );
  o21ai_0 U13653 ( .A1(n14527), .A2(n14528), .B1(n10749), .Y(n14515) );
  nand4_1 U13654 ( .A(n14471), .B(n14328), .C(n14481), .D(n14529), .Y(n14528)
         );
  and3_1 U13655 ( .A(n14530), .B(n10761), .C(n14347), .X(n14529) );
  inv_1 U13656 ( .A(n14531), .Y(n14347) );
  a21oi_1 U13657 ( .A1(n14532), .A2(n14533), .B1(n14534), .Y(n14328) );
  inv_1 U13658 ( .A(n14535), .Y(n14471) );
  o21ai_0 U13659 ( .A1(n14536), .A2(n14473), .B1(n14537), .Y(n14535) );
  nand4_1 U13660 ( .A(n14538), .B(n14395), .C(n14336), .D(n14539), .Y(n14527)
         );
  nor3_1 U13661 ( .A(n14540), .B(n14541), .C(n14299), .Y(n14539) );
  inv_1 U13662 ( .A(n14446), .Y(n14299) );
  nor4_1 U13663 ( .A(n14542), .B(n14543), .C(n14544), .D(n14545), .Y(n14514)
         );
  inv_1 U13664 ( .A(n14546), .Y(n14544) );
  nand3_1 U13665 ( .A(n14327), .B(n14293), .C(n14456), .Y(n14543) );
  and3_1 U13666 ( .A(n14319), .B(n14484), .C(n14375), .X(n14456) );
  and2_0 U13667 ( .A(n14547), .B(n14548), .X(n14327) );
  nand4_1 U13668 ( .A(n14320), .B(n10758), .C(n14486), .D(n14549), .Y(n14542)
         );
  nor2_1 U13669 ( .A(n10755), .B(n14550), .Y(n14549) );
  o211ai_1 U13670 ( .A1(n14551), .A2(n12842), .B1(n14400), .C1(n14552), .Y(
        n10379) );
  mux2i_1 U13671 ( .A0(n12847), .A1(n14553), .S(n14554), .Y(n14552) );
  nor4_1 U13672 ( .A(n14555), .B(n10769), .C(n14436), .D(n14545), .Y(n14554)
         );
  nand3_1 U13673 ( .A(n14332), .B(n14368), .C(n14445), .Y(n14545) );
  nand4_1 U13674 ( .A(n14334), .B(n14537), .C(n14470), .D(n14354), .Y(n14436)
         );
  nand4_1 U13675 ( .A(n14556), .B(n14344), .C(n14375), .D(n14557), .Y(n10769)
         );
  nor4_1 U13676 ( .A(n14558), .B(n14490), .C(n14491), .D(n14559), .Y(n14557)
         );
  inv_1 U13677 ( .A(n14395), .Y(n14558) );
  and3_1 U13678 ( .A(n14513), .B(n14306), .C(n14560), .X(n14344) );
  nand2_1 U13679 ( .A(n14561), .B(n14562), .Y(n14306) );
  inv_1 U13680 ( .A(n14283), .Y(n14556) );
  nand2_1 U13681 ( .A(n14510), .B(n14563), .Y(n14283) );
  and4_1 U13682 ( .A(n14564), .B(n14551), .C(n14565), .D(n10766), .X(n14553)
         );
  nand4_1 U13683 ( .A(n14566), .B(n14346), .C(n14567), .D(n14568), .Y(n10766)
         );
  nor4_1 U13684 ( .A(n14569), .B(n14444), .C(n14386), .D(n14409), .Y(n14568)
         );
  nand4_1 U13685 ( .A(n14320), .B(n14336), .C(n14570), .D(n14571), .Y(n14386)
         );
  and4_1 U13686 ( .A(n14572), .B(n14560), .C(n14314), .D(n14279), .X(n14571)
         );
  a211oi_1 U13687 ( .A1(n14573), .A2(n14574), .B1(n14575), .C1(n14491), .Y(
        n14279) );
  a21oi_1 U13688 ( .A1(n14576), .A2(n14574), .B1(n14526), .Y(n14314) );
  nor2_1 U13689 ( .A(n14349), .B(n14577), .Y(n14526) );
  a211oi_1 U13690 ( .A1(n14578), .A2(n14579), .B1(n14450), .C1(n12850), .Y(
        n14560) );
  inv_1 U13691 ( .A(n14465), .Y(n12850) );
  nand3_1 U13692 ( .A(n14580), .B(n14578), .C(n14581), .Y(n14465) );
  nor3_1 U13693 ( .A(n14536), .B(n14577), .C(n12848), .Y(n14450) );
  nor3_1 U13694 ( .A(n14490), .B(n14288), .C(n14289), .Y(n14570) );
  inv_1 U13695 ( .A(n14521), .Y(n14289) );
  nand3_1 U13696 ( .A(n14582), .B(n14578), .C(n14583), .Y(n14521) );
  inv_1 U13697 ( .A(n14498), .Y(n14490) );
  nand3_1 U13698 ( .A(n14584), .B(n14585), .C(n14586), .Y(n14320) );
  nand3_1 U13699 ( .A(n14530), .B(n14587), .C(n14345), .Y(n14569) );
  nor2_1 U13700 ( .A(n10768), .B(n14454), .Y(n14345) );
  inv_1 U13701 ( .A(n14388), .Y(n14454) );
  nand3_1 U13702 ( .A(n14586), .B(n14588), .C(n14589), .Y(n14388) );
  inv_1 U13703 ( .A(n14411), .Y(n10768) );
  nand3_1 U13704 ( .A(n14590), .B(n14578), .C(n14584), .Y(n14411) );
  inv_1 U13705 ( .A(n14414), .Y(n14587) );
  nand3_1 U13706 ( .A(n14358), .B(n14440), .C(n14319), .Y(n14414) );
  nand3_1 U13707 ( .A(n14591), .B(n14592), .C(n14593), .Y(n14319) );
  and4_1 U13708 ( .A(n14302), .B(n14594), .C(n14321), .D(n14595), .X(n14530)
         );
  and2_0 U13709 ( .A(n14423), .B(n14387), .X(n14595) );
  and4_1 U13710 ( .A(n14513), .B(n14467), .C(n10765), .D(n14416), .X(n14387)
         );
  nand3_1 U13711 ( .A(n14596), .B(n14597), .C(n14598), .Y(n14513) );
  nor2_1 U13712 ( .A(n14380), .B(n10767), .Y(n14423) );
  inv_1 U13713 ( .A(n14353), .Y(n10767) );
  nand2_1 U13714 ( .A(n14599), .B(n14580), .Y(n14353) );
  inv_1 U13715 ( .A(n14600), .Y(n14380) );
  nand3_1 U13716 ( .A(n14593), .B(n14573), .C(n14601), .Y(n14321) );
  nor3_1 U13717 ( .A(n14379), .B(n14477), .C(n14489), .Y(n14567) );
  inv_1 U13718 ( .A(n10758), .Y(n14489) );
  inv_1 U13719 ( .A(n14510), .Y(n14477) );
  inv_1 U13720 ( .A(n14363), .Y(n14379) );
  nand3_1 U13721 ( .A(n14585), .B(n14580), .C(n14602), .Y(n14363) );
  nor2_1 U13722 ( .A(n14418), .B(n14381), .Y(n14346) );
  inv_1 U13723 ( .A(n14603), .Y(n14418) );
  nor2_1 U13724 ( .A(n14503), .B(n14559), .Y(n14566) );
  nand4_1 U13725 ( .A(n14303), .B(n14301), .C(n14474), .D(n14604), .Y(n14559)
         );
  nor2_1 U13726 ( .A(n14531), .B(n14282), .Y(n14604) );
  nand4_1 U13727 ( .A(n14548), .B(n14424), .C(n14364), .D(n14438), .Y(n14282)
         );
  nand2_1 U13728 ( .A(n14394), .B(n14317), .Y(n14531) );
  nand3_1 U13729 ( .A(n14605), .B(n14597), .C(n14606), .Y(n14317) );
  nor4_1 U13730 ( .A(n12851), .B(n14449), .C(n14453), .D(n14501), .Y(n14474)
         );
  inv_1 U13731 ( .A(n14415), .Y(n14449) );
  inv_1 U13732 ( .A(n14447), .Y(n12851) );
  nand2_1 U13733 ( .A(n14607), .B(n14590), .Y(n14447) );
  nand2_1 U13734 ( .A(n14574), .B(n14585), .Y(n14303) );
  nand4_1 U13735 ( .A(n14313), .B(n14435), .C(n14538), .D(n14354), .Y(n14503)
         );
  nand3_1 U13736 ( .A(n14583), .B(n14608), .C(n14609), .Y(n14354) );
  and3_1 U13737 ( .A(n14425), .B(n14359), .C(n14331), .X(n14435) );
  and4_1 U13738 ( .A(n14352), .B(n14332), .C(n14294), .D(n14610), .X(n14425)
         );
  and3_1 U13739 ( .A(n14284), .B(n14547), .C(n14307), .X(n14610) );
  nand3_1 U13740 ( .A(n14611), .B(n14612), .C(n14609), .Y(n14307) );
  inv_1 U13741 ( .A(n14534), .Y(n14294) );
  nand3_1 U13742 ( .A(n14613), .B(n14614), .C(n14565), .Y(n14534) );
  and3_1 U13743 ( .A(n14333), .B(n10697), .C(n14441), .X(n14564) );
  inv_1 U13744 ( .A(n10747), .Y(n12847) );
  and4_1 U13745 ( .A(n14615), .B(n14329), .C(n14481), .D(n14616), .X(n14551)
         );
  nor4_1 U13746 ( .A(n14617), .B(n14618), .C(n10754), .D(n10755), .Y(n14616)
         );
  nand4_1 U13747 ( .A(n14350), .B(n14316), .C(n14351), .D(n14619), .Y(n10755)
         );
  nand3_1 U13748 ( .A(n14605), .B(n14298), .C(n14593), .Y(n14350) );
  nand4_1 U13749 ( .A(n14277), .B(n14467), .C(n14308), .D(n14416), .Y(n10754)
         );
  nand3_1 U13750 ( .A(n14620), .B(n14621), .C(n14611), .Y(n14308) );
  and4_1 U13751 ( .A(n14483), .B(n14507), .C(n14603), .D(n14336), .X(n14277)
         );
  nand3_1 U13752 ( .A(n14588), .B(n14576), .C(n14622), .Y(n14507) );
  inv_1 U13753 ( .A(n14623), .Y(n14483) );
  o21ai_0 U13754 ( .A1(n14455), .A2(n14361), .B1(n14367), .Y(n14623) );
  nand3_1 U13755 ( .A(n14586), .B(n14590), .C(n14601), .Y(n14367) );
  nor3_1 U13756 ( .A(n14624), .B(n14625), .C(n14626), .Y(n14618) );
  inv_1 U13757 ( .A(n14352), .Y(n14617) );
  nand2_1 U13758 ( .A(n14627), .B(n14628), .Y(n14352) );
  nor2_1 U13759 ( .A(n14629), .B(n14630), .Y(n14329) );
  inv_1 U13760 ( .A(n14406), .Y(n14615) );
  nand4_1 U13761 ( .A(n10759), .B(n10765), .C(n10761), .D(n14631), .Y(n14406)
         );
  nor2_1 U13762 ( .A(n10764), .B(n14437), .Y(n14631) );
  nand4_1 U13763 ( .A(n14362), .B(n14302), .C(n14366), .D(n14389), .Y(n14437)
         );
  nand4_1 U13764 ( .A(n14632), .B(n14286), .C(n14446), .D(n14594), .Y(n10764)
         );
  nand2_1 U13765 ( .A(n14633), .B(n14593), .Y(n14594) );
  o21ai_0 U13766 ( .A1(n14633), .A2(n14634), .B1(n14586), .Y(n14286) );
  nor2_1 U13767 ( .A(n10756), .B(n12848), .Y(n14634) );
  and2_0 U13768 ( .A(n14589), .B(n14582), .X(n14633) );
  nand2_1 U13769 ( .A(n14601), .B(n14599), .Y(n14632) );
  a21oi_1 U13770 ( .A1(n14635), .A2(n14636), .B1(n14512), .Y(n10761) );
  and3_1 U13771 ( .A(n14578), .B(n14573), .C(n14580), .X(n14512) );
  nand2_1 U13772 ( .A(n14298), .B(n14637), .Y(n10765) );
  a21oi_1 U13773 ( .A1(n14597), .A2(n14638), .B1(n14540), .Y(n10759) );
  inv_1 U13774 ( .A(n14278), .Y(n14540) );
  nand3_1 U13775 ( .A(n14582), .B(n14578), .C(n14585), .Y(n14278) );
  nor2_1 U13776 ( .A(n14455), .B(n14577), .Y(n14638) );
  o221ai_1 U13777 ( .A1(n14639), .A2(n10747), .B1(n14640), .B2(n12842), .C1(
        n14641), .Y(n10378) );
  a21oi_1 U13778 ( .A1(n10697), .A2(n14642), .B1(n14643), .Y(n14641) );
  inv_1 U13779 ( .A(n14400), .Y(n14643) );
  nand3_1 U13780 ( .A(n14601), .B(n14644), .C(n10749), .Y(n14400) );
  inv_1 U13781 ( .A(n12842), .Y(n10749) );
  inv_1 U13782 ( .A(n12848), .Y(n14601) );
  nand4_1 U13783 ( .A(n24042), .B(n12472), .C(n12355), .D(n12316), .Y(n12848)
         );
  nand4_1 U13784 ( .A(n14645), .B(n14375), .C(n14646), .D(n14647), .Y(n14642)
         );
  nor4_1 U13785 ( .A(n14648), .B(n14555), .C(n14491), .D(n14649), .Y(n14647)
         );
  inv_1 U13786 ( .A(n14438), .Y(n14649) );
  nand3_1 U13787 ( .A(n14602), .B(n14650), .C(n14598), .Y(n14438) );
  nor3_1 U13788 ( .A(n14651), .B(n14652), .C(n14653), .Y(n14491) );
  inv_1 U13789 ( .A(n14284), .Y(n14555) );
  nand2_1 U13790 ( .A(n14627), .B(n14612), .Y(n14284) );
  nand3_1 U13791 ( .A(n14600), .B(n14547), .C(n14498), .Y(n14648) );
  nand3_1 U13792 ( .A(n14620), .B(n14621), .C(n14654), .Y(n14498) );
  nand3_1 U13793 ( .A(n14611), .B(n14612), .C(n14655), .Y(n14547) );
  nand2_1 U13794 ( .A(n14644), .B(n14591), .Y(n14600) );
  inv_1 U13795 ( .A(n14455), .Y(n14591) );
  nand3_1 U13796 ( .A(n12355), .B(n14656), .C(n14657), .Y(n14455) );
  nor3_1 U13797 ( .A(n14463), .B(n14300), .C(n14396), .Y(n14646) );
  nand3_1 U13798 ( .A(n14358), .B(n14510), .C(n14351), .Y(n14396) );
  nand3_1 U13799 ( .A(n14657), .B(n14658), .C(n14659), .Y(n14351) );
  nand3_1 U13800 ( .A(n14636), .B(n14660), .C(n14598), .Y(n14510) );
  and3_1 U13801 ( .A(n14657), .B(n14658), .C(n14661), .X(n14598) );
  nand2_1 U13802 ( .A(n14662), .B(n14611), .Y(n14358) );
  nand3_1 U13803 ( .A(n14538), .B(n14416), .C(n14467), .Y(n14300) );
  nand2_1 U13804 ( .A(n14297), .B(n14620), .Y(n14467) );
  nand2_1 U13805 ( .A(n14562), .B(n14659), .Y(n14416) );
  inv_1 U13806 ( .A(n14629), .Y(n14538) );
  nor3_1 U13807 ( .A(n14626), .B(n14663), .C(n14624), .Y(n14629) );
  nand2_1 U13808 ( .A(n14546), .B(n14563), .Y(n14463) );
  nand2_1 U13809 ( .A(n14561), .B(n14664), .Y(n14563) );
  nor3_1 U13810 ( .A(n14665), .B(n14652), .C(n14666), .Y(n14561) );
  a21oi_1 U13811 ( .A1(n14576), .A2(n14574), .B1(n14667), .Y(n14546) );
  inv_1 U13812 ( .A(n14440), .Y(n14667) );
  nand2_1 U13813 ( .A(n14579), .B(n14586), .Y(n14440) );
  inv_1 U13814 ( .A(n14473), .Y(n14579) );
  a21oi_1 U13815 ( .A1(n14298), .A2(n14297), .B1(n14668), .Y(n14375) );
  inv_1 U13816 ( .A(n14360), .Y(n14668) );
  nand4_1 U13817 ( .A(n14620), .B(n14661), .C(n14636), .D(n14660), .Y(n14360)
         );
  and2_0 U13818 ( .A(n14614), .B(n14313), .X(n14645) );
  and4_1 U13819 ( .A(n14334), .B(n14537), .C(n14366), .D(n14669), .X(n14313)
         );
  nor3_1 U13820 ( .A(n14385), .B(n14630), .C(n14550), .Y(n14669) );
  nand4_1 U13821 ( .A(n14441), .B(n14470), .C(n14333), .D(n14389), .Y(n14550)
         );
  nand3_1 U13822 ( .A(n14654), .B(n14670), .C(n14655), .Y(n14389) );
  nand3_1 U13823 ( .A(n14532), .B(n14671), .C(n14655), .Y(n14333) );
  nand3_1 U13824 ( .A(n14576), .B(n14670), .C(n14609), .Y(n14470) );
  nand3_1 U13825 ( .A(n14611), .B(n14628), .C(n14655), .Y(n14441) );
  nor3_1 U13826 ( .A(n14672), .B(n14673), .C(n14624), .Y(n14630) );
  o21ai_0 U13827 ( .A1(n14653), .A2(n14674), .B1(n14368), .Y(n14385) );
  nand2_1 U13828 ( .A(n14533), .B(n14605), .Y(n14368) );
  nand2_1 U13829 ( .A(n14533), .B(n14583), .Y(n14366) );
  nand3_1 U13830 ( .A(n14589), .B(n14671), .C(n14655), .Y(n14537) );
  nand3_1 U13831 ( .A(n14589), .B(n14608), .C(n14609), .Y(n14334) );
  nand3_1 U13832 ( .A(n14675), .B(n14676), .C(n14627), .Y(n14614) );
  and2_0 U13833 ( .A(n14655), .B(n14581), .X(n14627) );
  nand2_1 U13834 ( .A(n14677), .B(n10697), .Y(n12842) );
  nor4_1 U13835 ( .A(n14678), .B(n14679), .C(n14499), .D(n14680), .Y(n14640)
         );
  inv_1 U13836 ( .A(n14481), .Y(n14680) );
  a21oi_1 U13837 ( .A1(n14585), .A2(n14607), .B1(n14281), .Y(n14481) );
  o32ai_1 U13838 ( .A1(n14681), .A2(n14577), .A3(n14536), .B1(n14348), .B2(
        n10757), .Y(n14281) );
  inv_1 U13839 ( .A(n10757), .Y(n14607) );
  inv_1 U13840 ( .A(n10756), .Y(n14585) );
  nand2_1 U13841 ( .A(n14682), .B(n14683), .Y(n10756) );
  nand2_1 U13842 ( .A(n14302), .B(n10758), .Y(n14499) );
  nand3_1 U13843 ( .A(n14592), .B(n14636), .C(n14588), .Y(n10758) );
  nand3_1 U13844 ( .A(n14293), .B(n14572), .C(n14315), .Y(n14679) );
  inv_1 U13845 ( .A(n14357), .Y(n14315) );
  nand2_1 U13846 ( .A(n14445), .B(n14395), .Y(n14357) );
  nand2_1 U13847 ( .A(n14297), .B(n14664), .Y(n14395) );
  and2_0 U13848 ( .A(n14684), .B(n14602), .X(n14297) );
  nand3_1 U13849 ( .A(n14684), .B(n14597), .C(n14606), .Y(n14445) );
  and2_0 U13850 ( .A(n10771), .B(n14484), .X(n14572) );
  nand2_1 U13851 ( .A(n14644), .B(n14582), .Y(n14484) );
  nand2_1 U13852 ( .A(n14593), .B(n14635), .Y(n10771) );
  inv_1 U13853 ( .A(n14444), .Y(n14293) );
  o21ai_0 U13854 ( .A1(n10757), .A2(n14672), .B1(n14422), .Y(n14444) );
  nand3_1 U13855 ( .A(n14588), .B(n14576), .C(n14597), .Y(n14422) );
  inv_1 U13856 ( .A(n14589), .Y(n14672) );
  nand2_1 U13857 ( .A(n14588), .B(n14578), .Y(n10757) );
  inv_1 U13858 ( .A(n14472), .Y(n14578) );
  nand2_1 U13859 ( .A(n14670), .B(n14685), .Y(n14472) );
  nand4_1 U13860 ( .A(n14548), .B(n14424), .C(n14394), .D(n14686), .Y(n14678)
         );
  nor3_1 U13861 ( .A(n14392), .B(n14453), .C(n14381), .Y(n14686) );
  inv_1 U13862 ( .A(n14524), .Y(n14381) );
  nand2_1 U13863 ( .A(n14584), .B(n14599), .Y(n14524) );
  inv_1 U13864 ( .A(n14361), .Y(n14599) );
  nand2_1 U13865 ( .A(n14590), .B(n14636), .Y(n14361) );
  inv_1 U13866 ( .A(n14305), .Y(n14453) );
  nand2_1 U13867 ( .A(n14562), .B(n14637), .Y(n14305) );
  and3_1 U13868 ( .A(n12472), .B(n12355), .C(n14657), .X(n14562) );
  inv_1 U13869 ( .A(n14301), .Y(n14392) );
  nand3_1 U13870 ( .A(n14298), .B(n14602), .C(n14605), .Y(n14301) );
  nand3_1 U13871 ( .A(n14593), .B(n14298), .C(n14684), .Y(n14394) );
  nor2_1 U13872 ( .A(n14666), .B(n14687), .Y(n14684) );
  nand3_1 U13873 ( .A(n14620), .B(n14597), .C(n14532), .Y(n14424) );
  nand4_1 U13874 ( .A(n14606), .B(n14661), .C(n14622), .D(n14682), .Y(n14548)
         );
  nand2_1 U13875 ( .A(inData[21]), .B(n10697), .Y(n10747) );
  nor4_1 U13876 ( .A(n14688), .B(n14689), .C(n14409), .D(n14485), .Y(n14639)
         );
  nand4_1 U13877 ( .A(n14613), .B(n14332), .C(n14565), .D(n14690), .Y(n14485)
         );
  nor3_1 U13878 ( .A(n14541), .B(n14288), .C(n14575), .Y(n14690) );
  inv_1 U13879 ( .A(n10773), .Y(n14575) );
  nand2_1 U13880 ( .A(n14581), .B(n14574), .Y(n10773) );
  inv_1 U13881 ( .A(n14349), .Y(n14574) );
  nand2_1 U13882 ( .A(n14593), .B(n14588), .Y(n14349) );
  nor4_1 U13883 ( .A(n14656), .B(n14691), .C(n14692), .D(n24042), .Y(n14588)
         );
  inv_1 U13884 ( .A(n14619), .Y(n14288) );
  nand2_1 U13885 ( .A(n14659), .B(n14664), .Y(n14619) );
  and3_1 U13886 ( .A(n12472), .B(n14691), .C(n14657), .X(n14664) );
  nor2_1 U13887 ( .A(n14693), .B(n12316), .Y(n14657) );
  and3_1 U13888 ( .A(n14621), .B(n14650), .C(n14661), .X(n14659) );
  inv_1 U13889 ( .A(n14364), .Y(n14541) );
  nand3_1 U13890 ( .A(n14654), .B(n14586), .C(n14606), .Y(n14364) );
  nand3_1 U13891 ( .A(n14581), .B(n14628), .C(n14609), .Y(n14565) );
  inv_1 U13892 ( .A(n14694), .Y(n14628) );
  nand3_1 U13893 ( .A(n14532), .B(n14671), .C(n14609), .Y(n14332) );
  nand3_1 U13894 ( .A(n14654), .B(n14670), .C(n14609), .Y(n14613) );
  inv_1 U13895 ( .A(n14695), .Y(n14670) );
  o211ai_1 U13896 ( .A1(n14536), .A2(n14473), .B1(n10772), .C1(n14378), .Y(
        n14409) );
  nand3_1 U13897 ( .A(n14592), .B(n14580), .C(n14622), .Y(n14378) );
  inv_1 U13898 ( .A(n14577), .Y(n14592) );
  nand2_1 U13899 ( .A(n14650), .B(n14683), .Y(n14577) );
  nand3_1 U13900 ( .A(n14584), .B(n14573), .C(n14593), .Y(n10772) );
  nor3_1 U13901 ( .A(n24045), .B(n24046), .C(n14696), .Y(n14593) );
  inv_1 U13902 ( .A(n14348), .Y(n14573) );
  nand2_1 U13903 ( .A(n14683), .B(n14660), .Y(n14348) );
  inv_1 U13904 ( .A(n14681), .Y(n14584) );
  nand3_1 U13905 ( .A(n12316), .B(n14658), .C(n24042), .Y(n14681) );
  nand2_1 U13906 ( .A(n14583), .B(n14580), .Y(n14473) );
  nor2_1 U13907 ( .A(n14687), .B(n14697), .Y(n14583) );
  nand3_1 U13908 ( .A(n14316), .B(n14362), .C(n14331), .Y(n14689) );
  inv_1 U13909 ( .A(n14398), .Y(n14331) );
  nand2_1 U13910 ( .A(n14486), .B(n14285), .Y(n14398) );
  nand2_1 U13911 ( .A(n14662), .B(n14581), .Y(n14285) );
  nor3_1 U13912 ( .A(n14698), .B(n24047), .C(n14624), .Y(n14662) );
  nand2_1 U13913 ( .A(n14533), .B(n14589), .Y(n14486) );
  nor2_1 U13914 ( .A(n14665), .B(n14697), .Y(n14589) );
  inv_1 U13915 ( .A(n14674), .Y(n14533) );
  nand2_1 U13916 ( .A(n14655), .B(n14608), .Y(n14674) );
  inv_1 U13917 ( .A(n14699), .Y(n14608) );
  and3_1 U13918 ( .A(n12472), .B(n14691), .C(n14700), .X(n14655) );
  nand2_1 U13919 ( .A(n14620), .B(n14637), .Y(n14362) );
  nand3_1 U13920 ( .A(n14298), .B(n14586), .C(n14654), .Y(n14316) );
  nor2_1 U13921 ( .A(n14701), .B(n14702), .Y(n14654) );
  nand4_1 U13922 ( .A(n14415), .B(n14603), .C(n14446), .D(n14703), .Y(n14688)
         );
  nor3_1 U13923 ( .A(n14704), .B(n14523), .C(n14501), .Y(n14703) );
  and2_0 U13924 ( .A(n14644), .B(n14580), .X(n14501) );
  and3_1 U13925 ( .A(n14658), .B(n14693), .C(n12316), .X(n14580) );
  inv_1 U13926 ( .A(n12849), .Y(n14644) );
  nand2_1 U13927 ( .A(n14590), .B(n14622), .Y(n12849) );
  inv_1 U13928 ( .A(n14536), .Y(n14622) );
  nand2_1 U13929 ( .A(n14612), .B(n14685), .Y(n14536) );
  inv_1 U13930 ( .A(n14625), .Y(n14612) );
  nor2_1 U13931 ( .A(n14687), .B(n14705), .Y(n14590) );
  inv_1 U13932 ( .A(n14359), .Y(n14523) );
  nand2_1 U13933 ( .A(n14609), .B(n14706), .Y(n14359) );
  o22ai_1 U13934 ( .A1(n14625), .A2(n14626), .B1(n14699), .B2(n14653), .Y(
        n14706) );
  inv_1 U13935 ( .A(n14532), .Y(n14653) );
  nor2_1 U13936 ( .A(n14701), .B(n14665), .Y(n14532) );
  inv_1 U13937 ( .A(n14581), .Y(n14626) );
  nor2_1 U13938 ( .A(n14697), .B(n14707), .Y(n14581) );
  inv_1 U13939 ( .A(n14624), .Y(n14609) );
  nand3_1 U13940 ( .A(n12355), .B(n14656), .C(n14700), .Y(n14624) );
  nor3_1 U13941 ( .A(n14693), .B(n14692), .C(n14685), .Y(n14700) );
  inv_1 U13942 ( .A(n12316), .Y(n14692) );
  inv_1 U13943 ( .A(n14336), .Y(n14704) );
  nand2_1 U13944 ( .A(n14606), .B(n14637), .Y(n14336) );
  and3_1 U13945 ( .A(n14621), .B(n14660), .C(n14661), .X(n14637) );
  nor2_1 U13946 ( .A(n14699), .B(n24045), .Y(n14621) );
  nand4_1 U13947 ( .A(n14298), .B(n14586), .C(n14661), .D(n14650), .Y(n14446)
         );
  nor2_1 U13948 ( .A(n14694), .B(n24045), .Y(n14586) );
  inv_1 U13949 ( .A(n14651), .Y(n14298) );
  nand2_1 U13950 ( .A(n14708), .B(n14658), .Y(n14651) );
  nor2_1 U13951 ( .A(n12355), .B(n12472), .Y(n14658) );
  nand3_1 U13952 ( .A(n14620), .B(n14602), .C(n14605), .Y(n14603) );
  nor2_1 U13953 ( .A(n14701), .B(n14687), .Y(n14605) );
  nor2_1 U13954 ( .A(n14663), .B(n24045), .Y(n14602) );
  and3_1 U13955 ( .A(n12355), .B(n14708), .C(n12472), .X(n14620) );
  nand2_1 U13956 ( .A(n14597), .B(n14635), .Y(n14415) );
  and2_0 U13957 ( .A(n14576), .B(n14582), .X(n14635) );
  and3_1 U13958 ( .A(n14708), .B(n14656), .C(n12355), .X(n14582) );
  inv_1 U13959 ( .A(n12472), .Y(n14656) );
  nor2_1 U13960 ( .A(n14702), .B(n14697), .Y(n14576) );
  inv_1 U13961 ( .A(n14652), .Y(n14597) );
  nand3_1 U13962 ( .A(n14685), .B(n14676), .C(n14675), .Y(n14652) );
  o221ai_1 U13963 ( .A1(n14709), .A2(n14710), .B1(n14711), .B2(n10977), .C1(
        n14712), .Y(n10377) );
  a21oi_1 U13964 ( .A1(n14302), .A2(n14713), .B1(n14714), .Y(n14712) );
  nand4_1 U13965 ( .A(n14715), .B(n14716), .C(n14717), .D(n14718), .Y(n14713)
         );
  nor4_1 U13966 ( .A(n14719), .B(n14720), .C(n14721), .D(n14722), .Y(n14718)
         );
  nand3_1 U13967 ( .A(n14723), .B(n14724), .C(n14725), .Y(n14719) );
  and3_1 U13968 ( .A(n14726), .B(n14727), .C(n14728), .X(n14717) );
  inv_1 U13969 ( .A(n14729), .Y(n14715) );
  nor4_1 U13970 ( .A(n14730), .B(n14731), .C(n14732), .D(n14733), .Y(n14711)
         );
  nand3_1 U13971 ( .A(n11030), .B(n14734), .C(n14735), .Y(n14731) );
  nand4_1 U13972 ( .A(n14736), .B(n14737), .C(n14738), .D(n14739), .Y(n14730)
         );
  and3_1 U13973 ( .A(n11024), .B(n14740), .C(n14741), .X(n14739) );
  nor4_1 U13974 ( .A(n14742), .B(n14743), .C(n11027), .D(n14744), .Y(n14709)
         );
  nand4_1 U13975 ( .A(n14745), .B(n14746), .C(n14747), .D(n14748), .Y(n11027)
         );
  nor3_1 U13976 ( .A(n14749), .B(n14750), .C(n14751), .Y(n14748) );
  nand3_1 U13977 ( .A(n14752), .B(n14753), .C(n14754), .Y(n14749) );
  nor3_1 U13978 ( .A(n14755), .B(n14756), .C(n14757), .Y(n14747) );
  inv_1 U13979 ( .A(n14758), .Y(n14756) );
  inv_1 U13980 ( .A(n14759), .Y(n14745) );
  nand2_1 U13981 ( .A(n14760), .B(n14761), .Y(n14743) );
  nand4_1 U13982 ( .A(n14762), .B(n14763), .C(n14764), .D(n14765), .Y(n14742)
         );
  nand4_1 U13983 ( .A(n14766), .B(n14767), .C(n14768), .D(n14769), .Y(n10376)
         );
  nand2_1 U13984 ( .A(n14770), .B(n14302), .Y(n14767) );
  nand4_1 U13985 ( .A(n14771), .B(n14772), .C(n14773), .D(n14774), .Y(n14770)
         );
  nor3_1 U13986 ( .A(n14775), .B(n14776), .C(n14777), .Y(n14774) );
  nand3_1 U13987 ( .A(n14723), .B(n14778), .C(n14779), .Y(n14775) );
  a21oi_1 U13988 ( .A1(n14780), .A2(n14781), .B1(n14782), .Y(n14773) );
  inv_1 U13989 ( .A(n14783), .Y(n14772) );
  mux2i_1 U13990 ( .A0(n14784), .A1(n14785), .S(n14786), .Y(n14766) );
  nor4_1 U13991 ( .A(n14787), .B(n14788), .C(n11029), .D(n14789), .Y(n14786)
         );
  nand3_1 U13992 ( .A(n14790), .B(n14736), .C(n14791), .Y(n14787) );
  nor4_1 U13993 ( .A(n14792), .B(n14793), .C(n14755), .D(n10998), .Y(n14785)
         );
  inv_1 U13994 ( .A(n14794), .Y(n14755) );
  nand2_1 U13995 ( .A(n14752), .B(n11006), .Y(n14793) );
  or4_1 U13996 ( .A(n14795), .B(n14796), .C(n14797), .D(n14710), .X(n14792) );
  o211ai_1 U13997 ( .A1(n14798), .A2(n10977), .B1(n14768), .C1(n14799), .Y(
        n10375) );
  mux2i_1 U13998 ( .A0(n10980), .A1(n14800), .S(n14801), .Y(n14799) );
  nor4_1 U13999 ( .A(n14802), .B(n14803), .C(n14804), .D(n14805), .Y(n14801)
         );
  nand3_1 U14000 ( .A(n14806), .B(n14807), .C(n14808), .Y(n14803) );
  nand4_1 U14001 ( .A(n14725), .B(n14809), .C(n14810), .D(n14754), .Y(n14802)
         );
  nor2_1 U14002 ( .A(n14811), .B(n14812), .Y(n14810) );
  nor4_1 U14003 ( .A(n14813), .B(n14814), .C(n10998), .D(n14815), .Y(n14800)
         );
  nand2_1 U14004 ( .A(n14816), .B(n14817), .Y(n14815) );
  nand3_1 U14005 ( .A(n14818), .B(n14798), .C(n14819), .Y(n14814) );
  inv_1 U14006 ( .A(n14820), .Y(n14819) );
  nand4_1 U14007 ( .A(n14821), .B(n14302), .C(n14791), .D(n14822), .Y(n14813)
         );
  nor3_1 U14008 ( .A(n14823), .B(n14824), .C(n14825), .Y(n14822) );
  and4_1 U14009 ( .A(n14826), .B(n14827), .C(n14828), .D(n14829), .X(n14798)
         );
  nor3_1 U14010 ( .A(n14830), .B(n14831), .C(n14832), .Y(n14829) );
  nand3_1 U14011 ( .A(n14737), .B(n14833), .C(n11003), .Y(n14830) );
  and3_1 U14012 ( .A(n14834), .B(n14835), .C(n10994), .X(n14828) );
  inv_1 U14013 ( .A(n14788), .Y(n14827) );
  nand3_1 U14014 ( .A(n14836), .B(n14837), .C(n14838), .Y(n14788) );
  nand4_1 U14015 ( .A(n14839), .B(n14840), .C(n14841), .D(n14842), .Y(n10374)
         );
  nor4_1 U14016 ( .A(n14843), .B(n14844), .C(n14845), .D(n14846), .Y(n14842)
         );
  o22ai_1 U14017 ( .A1(n14847), .A2(n14848), .B1(n14849), .B2(n14850), .Y(
        n14844) );
  a21oi_1 U14018 ( .A1(n14851), .A2(n14852), .B1(n14853), .Y(n14849) );
  a21oi_1 U14019 ( .A1(n14854), .A2(n14855), .B1(n14856), .Y(n14847) );
  inv_1 U14020 ( .A(n14857), .Y(n14854) );
  o221ai_1 U14021 ( .A1(n14858), .A2(n12466), .B1(n14859), .B2(n14860), .C1(
        n14861), .Y(n14843) );
  o21ai_0 U14022 ( .A1(n14862), .A2(n14863), .B1(n14864), .Y(n14861) );
  nor3_1 U14023 ( .A(n14865), .B(n14866), .C(n14867), .Y(n14860) );
  nand4_1 U14024 ( .A(n14868), .B(n14869), .C(n14870), .D(n14871), .Y(n14867)
         );
  nand3_1 U14025 ( .A(n14872), .B(n14873), .C(n14874), .Y(n14869) );
  nand3_1 U14026 ( .A(n14875), .B(n14876), .C(n14877), .Y(n14868) );
  nand4_1 U14027 ( .A(n14878), .B(n14879), .C(n14880), .D(n14881), .Y(n14866)
         );
  nand4_1 U14028 ( .A(n14882), .B(n14883), .C(n14884), .D(n14885), .Y(n14865)
         );
  nor3_1 U14029 ( .A(n14886), .B(n14887), .C(n14888), .Y(n14885) );
  o22ai_1 U14030 ( .A1(n14889), .A2(n14857), .B1(n14890), .B2(n14891), .Y(
        n14886) );
  inv_1 U14031 ( .A(n14892), .Y(n14883) );
  inv_1 U14032 ( .A(n14893), .Y(n14841) );
  o221ai_1 U14033 ( .A1(n14894), .A2(n14895), .B1(n14896), .B2(n14897), .C1(
        n14898), .Y(n14893) );
  nor2_1 U14034 ( .A(n14899), .B(n14900), .Y(n14839) );
  inv_1 U14035 ( .A(n14901), .Y(n14899) );
  nand4_1 U14036 ( .A(n14902), .B(n14903), .C(n14904), .D(n14905), .Y(n10373)
         );
  nor3_1 U14037 ( .A(n14906), .B(n14845), .C(n14907), .Y(n14905) );
  and4_1 U14038 ( .A(n14908), .B(n14852), .C(n14909), .D(n24036), .X(n14845)
         );
  o32ai_1 U14039 ( .A1(n14857), .A2(n12466), .A3(n14889), .B1(n14859), .B2(
        n14910), .Y(n14906) );
  nor4_1 U14040 ( .A(n14911), .B(n14912), .C(n14913), .D(n14914), .Y(n14910)
         );
  nand4_1 U14041 ( .A(n14915), .B(n14916), .C(n14917), .D(n14918), .Y(n14911)
         );
  nand4_1 U14042 ( .A(n14919), .B(n14920), .C(n23892), .D(n10774), .Y(n14916)
         );
  nand2_1 U14043 ( .A(n14921), .B(n23837), .Y(n14915) );
  a222oi_1 U14044 ( .A1(n14922), .A2(n14923), .B1(n14924), .B2(n14925), .C1(
        n14926), .C2(n14864), .Y(n14904) );
  nor3_1 U14045 ( .A(n14927), .B(n14928), .C(n14929), .Y(n14903) );
  nor3_1 U14046 ( .A(n14930), .B(n14931), .C(n14932), .Y(n14902) );
  nand4_1 U14047 ( .A(n14933), .B(n14934), .C(n14935), .D(n14936), .Y(n10372)
         );
  nor4_1 U14048 ( .A(n14937), .B(n14938), .C(n14939), .D(n14940), .Y(n14936)
         );
  inv_1 U14049 ( .A(n14941), .Y(n14939) );
  o211ai_1 U14050 ( .A1(n14942), .A2(n14943), .B1(n14898), .C1(n14944), .Y(
        n14938) );
  inv_1 U14051 ( .A(n14945), .Y(n14944) );
  a21oi_1 U14052 ( .A1(n14946), .A2(n14947), .B1(n14948), .Y(n14898) );
  or4_1 U14053 ( .A(n14949), .B(n14950), .C(n14951), .D(n14952), .X(n14937) );
  nor4_1 U14054 ( .A(n14953), .B(n14954), .C(n14955), .D(n14956), .Y(n14935)
         );
  inv_1 U14055 ( .A(n14957), .Y(n14953) );
  a21oi_1 U14056 ( .A1(n14958), .A2(n14924), .B1(n14959), .Y(n14957) );
  nor2_1 U14057 ( .A(n14960), .B(n14859), .Y(n14924) );
  o21ai_0 U14058 ( .A1(n14961), .A2(n23872), .B1(n14962), .Y(n14958) );
  a222oi_1 U14059 ( .A1(n14963), .A2(n14964), .B1(n14965), .B2(n14966), .C1(
        n14946), .C2(n14967), .Y(n14934) );
  o211ai_1 U14060 ( .A1(n14968), .A2(n14969), .B1(n14970), .C1(n14971), .Y(
        n14967) );
  inv_1 U14061 ( .A(n14972), .Y(n14971) );
  o21ai_0 U14062 ( .A1(n14973), .A2(n14962), .B1(n14974), .Y(n14966) );
  nand4_1 U14063 ( .A(n14975), .B(n14976), .C(n14977), .D(n14978), .Y(n14963)
         );
  nor2_1 U14064 ( .A(n14979), .B(n14980), .Y(n14978) );
  o32ai_1 U14065 ( .A1(n14981), .A2(n14982), .A3(n14983), .B1(n14984), .B2(
        n14973), .Y(n14980) );
  inv_1 U14066 ( .A(n14985), .Y(n14976) );
  a22oi_1 U14067 ( .A1(n14986), .A2(n14987), .B1(n12460), .B2(n14988), .Y(
        n14933) );
  nand4_1 U14068 ( .A(n14989), .B(n14990), .C(n14991), .D(n14992), .Y(n10371)
         );
  a211oi_1 U14069 ( .A1(n14993), .A2(n14864), .B1(n14994), .C1(n14995), .Y(
        n14992) );
  a21oi_1 U14070 ( .A1(n14996), .A2(n14879), .B1(n14997), .Y(n14995) );
  o22ai_1 U14071 ( .A1(n14850), .A2(n14998), .B1(n14859), .B2(n14999), .Y(
        n14994) );
  nor4_1 U14072 ( .A(n15000), .B(n15001), .C(n15002), .D(n15003), .Y(n14999)
         );
  o21ai_0 U14073 ( .A1(n14984), .A2(n14960), .B1(n14974), .Y(n15003) );
  and3_1 U14074 ( .A(n15004), .B(n14896), .C(n15005), .X(n14974) );
  a21oi_1 U14075 ( .A1(n14925), .A2(n14852), .B1(n15006), .Y(n15005) );
  o211ai_1 U14076 ( .A1(n15007), .A2(n15008), .B1(n15009), .C1(n15010), .Y(
        n15001) );
  nand4_1 U14077 ( .A(n15011), .B(n15012), .C(n15013), .D(n15014), .Y(n15000)
         );
  nor3_1 U14078 ( .A(n15015), .B(n15016), .C(n15017), .Y(n15014) );
  inv_1 U14079 ( .A(n15018), .Y(n15015) );
  inv_1 U14080 ( .A(n14878), .Y(n14993) );
  a222oi_1 U14081 ( .A1(n15019), .A2(n14908), .B1(n15020), .B2(n14922), .C1(
        n15021), .C2(n12460), .Y(n14991) );
  nor4_1 U14082 ( .A(n15022), .B(n14948), .C(n14927), .D(n14950), .Y(n14990)
         );
  o21ai_0 U14083 ( .A1(n14895), .A2(n15023), .B1(n15024), .Y(n14950) );
  nand3_1 U14084 ( .A(n15025), .B(n15026), .C(n15027), .Y(n14927) );
  a221oi_1 U14085 ( .A1(n15028), .A2(n14922), .B1(n14864), .B2(n15029), .C1(
        n14956), .Y(n15027) );
  nor2_1 U14086 ( .A(n15030), .B(n14897), .Y(n14956) );
  nand3_1 U14087 ( .A(n15031), .B(n15032), .C(n15033), .Y(n15029) );
  inv_1 U14088 ( .A(n15034), .Y(n15028) );
  inv_1 U14089 ( .A(n15035), .Y(n15026) );
  o211ai_1 U14090 ( .A1(n14997), .A2(n15036), .B1(n15037), .C1(n15038), .Y(
        n14948) );
  nor3_1 U14091 ( .A(n15039), .B(n15040), .C(n15041), .Y(n14989) );
  nand3_1 U14092 ( .A(n15042), .B(n15043), .C(n15044), .Y(n10370) );
  nor4_1 U14093 ( .A(n15045), .B(n15046), .C(n15047), .D(n15048), .Y(n15044)
         );
  a21oi_1 U14094 ( .A1(n15049), .A2(n15050), .B1(n12466), .Y(n15048) );
  a21oi_1 U14095 ( .A1(n15051), .A2(n14870), .B1(n14850), .Y(n15047) );
  o22ai_1 U14096 ( .A1(n14848), .A2(n15052), .B1(n14859), .B2(n15053), .Y(
        n15046) );
  nor4_1 U14097 ( .A(n15054), .B(n15055), .C(n15021), .D(n15056), .Y(n15053)
         );
  inv_1 U14098 ( .A(n14996), .Y(n15056) );
  nand3_1 U14099 ( .A(n15032), .B(n15057), .C(n15058), .Y(n15055) );
  or4_1 U14100 ( .A(n15059), .B(n15060), .C(n15061), .D(n14926), .X(n15054) );
  inv_1 U14101 ( .A(n15062), .Y(n14926) );
  nand3_1 U14102 ( .A(n15063), .B(n15037), .C(n15064), .Y(n15045) );
  nor3_1 U14103 ( .A(n15065), .B(n14955), .C(n15066), .Y(n15064) );
  or3_1 U14104 ( .A(n14897), .B(n15067), .C(n15068), .X(n15063) );
  nor3_1 U14105 ( .A(n15069), .B(n15035), .C(n15070), .Y(n15043) );
  o211ai_1 U14106 ( .A1(n12466), .A2(n15071), .B1(n15072), .C1(n15073), .Y(
        n15035) );
  inv_1 U14107 ( .A(n15074), .Y(n15072) );
  o22ai_1 U14108 ( .A1(n14997), .A2(n15075), .B1(n15076), .B2(n15077), .Y(
        n15069) );
  nor4_1 U14109 ( .A(n15040), .B(n15078), .C(n15079), .D(n15080), .Y(n15042)
         );
  nand2_1 U14110 ( .A(n15081), .B(n15082), .Y(n15040) );
  a221oi_1 U14111 ( .A1(n15083), .A2(n14908), .B1(n14946), .B2(n14972), .C1(
        n15084), .Y(n15082) );
  o211ai_1 U14112 ( .A1(n14982), .A2(n15085), .B1(n15086), .C1(n15087), .Y(
        n14972) );
  a222oi_1 U14113 ( .A1(n15088), .A2(n14964), .B1(n15089), .B2(n12460), .C1(
        n15090), .C2(n14922), .Y(n15081) );
  inv_1 U14114 ( .A(n15091), .Y(n15088) );
  nand4_1 U14115 ( .A(n15092), .B(n15093), .C(n15094), .D(n15095), .Y(n10369)
         );
  nor4_1 U14116 ( .A(n15096), .B(n15097), .C(n15098), .D(n15099), .Y(n15095)
         );
  inv_1 U14117 ( .A(n15100), .Y(n15099) );
  a221oi_1 U14118 ( .A1(n15101), .A2(n14946), .B1(n14947), .B2(n15102), .C1(
        n15103), .Y(n15094) );
  a21oi_1 U14119 ( .A1(n15104), .A2(n15105), .B1(n14859), .Y(n15103) );
  nor4_1 U14120 ( .A(n15106), .B(n14853), .C(n15107), .D(n14862), .Y(n15105)
         );
  inv_1 U14121 ( .A(n15031), .Y(n14862) );
  nand3_1 U14122 ( .A(n15009), .B(n15108), .C(n15071), .Y(n15106) );
  nor4_1 U14123 ( .A(n14979), .B(n15109), .C(n15110), .D(n15111), .Y(n15104)
         );
  o32ai_1 U14124 ( .A1(n15112), .A2(n14984), .A3(n15113), .B1(n14960), .B2(
        n15114), .Y(n15109) );
  nand2_1 U14125 ( .A(n15010), .B(n14996), .Y(n14979) );
  inv_1 U14126 ( .A(n14917), .Y(n14947) );
  inv_1 U14127 ( .A(n15087), .Y(n15101) );
  nor4_1 U14128 ( .A(n15115), .B(n14931), .C(n14949), .D(n15041), .Y(n15093)
         );
  o221ai_1 U14129 ( .A1(n15116), .A2(n15076), .B1(n14942), .B2(n15117), .C1(
        n15118), .Y(n15041) );
  inv_1 U14130 ( .A(n15119), .Y(n15118) );
  nor2_1 U14131 ( .A(n15120), .B(n14913), .Y(n15116) );
  nand2_1 U14132 ( .A(n15121), .B(n15122), .Y(n14913) );
  inv_1 U14133 ( .A(n14880), .Y(n15120) );
  nand3_1 U14134 ( .A(n15123), .B(n15124), .C(n15125), .Y(n14949) );
  nor4_1 U14135 ( .A(n15126), .B(n15127), .C(n15074), .D(n15128), .Y(n15125)
         );
  inv_1 U14136 ( .A(n15129), .Y(n15126) );
  a21oi_1 U14137 ( .A1(n14946), .A2(n15130), .B1(n15070), .Y(n15123) );
  o22ai_1 U14138 ( .A1(n14942), .A2(n15018), .B1(n14895), .B2(n15131), .Y(
        n15070) );
  or3_1 U14139 ( .A(n15132), .B(n15133), .C(n15134), .X(n14931) );
  a21oi_1 U14140 ( .A1(n15135), .A2(n14884), .B1(n14850), .Y(n15134) );
  inv_1 U14141 ( .A(n15136), .Y(n15133) );
  nor3_1 U14142 ( .A(n15137), .B(n15138), .C(n15139), .Y(n15092) );
  nand4_1 U14143 ( .A(n15140), .B(n15141), .C(n15142), .D(n15143), .Y(n10368)
         );
  nor4_1 U14144 ( .A(n15084), .B(n15144), .C(n15145), .D(n15146), .Y(n15143)
         );
  nor2_1 U14145 ( .A(n14859), .B(n15147), .Y(n15146) );
  nor3_1 U14146 ( .A(n15148), .B(n15060), .C(n15111), .Y(n15147) );
  nand2_1 U14147 ( .A(n15149), .B(n15150), .Y(n15111) );
  nand4_1 U14148 ( .A(n15151), .B(n15152), .C(n15153), .D(n15154), .Y(n15060)
         );
  and3_1 U14149 ( .A(n15155), .B(n14882), .C(n14975), .X(n15154) );
  inv_1 U14150 ( .A(n15156), .Y(n14975) );
  o211ai_1 U14151 ( .A1(n14889), .A2(n14857), .B1(n15117), .C1(n15033), .Y(
        n15156) );
  a21oi_1 U14152 ( .A1(n14852), .A2(n14925), .B1(n15020), .Y(n14882) );
  inv_1 U14153 ( .A(n15157), .Y(n15020) );
  a21oi_1 U14154 ( .A1(n14852), .A2(n15158), .B1(n15159), .Y(n15153) );
  o221ai_1 U14155 ( .A1(n14981), .A2(n15160), .B1(n14973), .B2(n14962), .C1(
        n15131), .Y(n15148) );
  nand2_1 U14156 ( .A(n15161), .B(n12462), .Y(n15160) );
  a21oi_1 U14157 ( .A1(n15162), .A2(n15163), .B1(n14848), .Y(n15145) );
  nor3_1 U14158 ( .A(n14960), .B(n14997), .C(n14962), .Y(n15084) );
  nor3_1 U14159 ( .A(n15164), .B(n15165), .C(n14928), .Y(n15142) );
  nand4_1 U14160 ( .A(n15166), .B(n15167), .C(n15168), .D(n15169), .Y(n14928)
         );
  a222oi_1 U14161 ( .A1(n15083), .A2(n14964), .B1(n15170), .B2(n15102), .C1(
        n15171), .C2(n12460), .Y(n15169) );
  inv_1 U14162 ( .A(n14998), .Y(n15171) );
  inv_1 U14163 ( .A(n15052), .Y(n15170) );
  inv_1 U14164 ( .A(n15172), .Y(n15083) );
  a22oi_1 U14165 ( .A1(n14908), .A2(n15173), .B1(n15174), .B2(n14965), .Y(
        n15168) );
  nand3_1 U14166 ( .A(n15075), .B(n14896), .C(n14996), .Y(n15173) );
  o21ai_0 U14167 ( .A1(n14850), .A2(n15077), .B1(n15175), .Y(n15164) );
  nor4_1 U14168 ( .A(n14952), .B(n15078), .C(n15176), .D(n15177), .Y(n15141)
         );
  or4_1 U14169 ( .A(n14954), .B(n15132), .C(n15128), .D(n15178), .X(n15078) );
  o32ai_1 U14170 ( .A1(n14973), .A2(n14997), .A3(n14984), .B1(n12466), .B2(
        n15179), .Y(n15178) );
  nor3_1 U14171 ( .A(n12466), .B(n15180), .C(n14857), .Y(n14954) );
  o221ai_1 U14172 ( .A1(n14848), .A2(n15050), .B1(n14942), .B2(n15091), .C1(
        n15181), .Y(n14952) );
  o21ai_0 U14173 ( .A1(n15182), .A2(n15183), .B1(n14964), .Y(n15181) );
  nand2_1 U14174 ( .A(n15031), .B(n15034), .Y(n15183) );
  nand4_1 U14175 ( .A(n23873), .B(n15184), .C(n15185), .D(n15186), .Y(n15031)
         );
  nor2_1 U14176 ( .A(n15187), .B(n15180), .Y(n15186) );
  nor3_1 U14177 ( .A(n15188), .B(n15189), .C(n15190), .Y(n15140) );
  nand4_1 U14178 ( .A(n15191), .B(n15192), .C(n15193), .D(n15194), .Y(n10367)
         );
  a221oi_1 U14179 ( .A1(n14965), .A2(n15002), .B1(n15195), .B2(n14964), .C1(
        n15196), .Y(n15194) );
  o211ai_1 U14180 ( .A1(n15197), .A2(n14895), .B1(n15198), .C1(n15199), .Y(
        n15196) );
  nand3_1 U14181 ( .A(n14855), .B(n15200), .C(n12460), .Y(n15198) );
  inv_1 U14182 ( .A(n15201), .Y(n15197) );
  o21ai_0 U14183 ( .A1(n15202), .A2(n15203), .B1(n15018), .Y(n15201) );
  nand3_1 U14184 ( .A(n14925), .B(n15204), .C(n15205), .Y(n15018) );
  nand4_1 U14185 ( .A(n15206), .B(n15049), .C(n15207), .D(n15208), .Y(n15195)
         );
  nor3_1 U14186 ( .A(n15209), .B(n14912), .C(n14923), .Y(n15208) );
  o221ai_1 U14187 ( .A1(n14984), .A2(n14973), .B1(n15067), .B2(n15068), .C1(
        n15210), .Y(n14912) );
  and3_1 U14188 ( .A(n15117), .B(n14870), .C(n15091), .X(n15210) );
  nand3_1 U14189 ( .A(n15211), .B(n15033), .C(n15212), .Y(n15209) );
  inv_1 U14190 ( .A(n14888), .Y(n15212) );
  nand3_1 U14191 ( .A(n15204), .B(n15213), .C(n15205), .Y(n15033) );
  nand3_1 U14192 ( .A(n15214), .B(n23895), .C(n15215), .Y(n15211) );
  and3_1 U14193 ( .A(n15004), .B(n15216), .C(n15075), .X(n15207) );
  o21ai_0 U14194 ( .A1(n14960), .A2(n15217), .B1(n15150), .Y(n15002) );
  a211oi_1 U14195 ( .A1(n15016), .A2(n15102), .B1(n15218), .C1(n15219), .Y(
        n15193) );
  o22ai_1 U14196 ( .A1(n14848), .A2(n15071), .B1(n14850), .B2(n15220), .Y(
        n15218) );
  nor4_1 U14197 ( .A(n15221), .B(n14932), .C(n15222), .D(n14900), .Y(n15192)
         );
  o211ai_1 U14198 ( .A1(n12466), .A2(n15058), .B1(n15223), .C1(n15224), .Y(
        n14900) );
  a211oi_1 U14199 ( .A1(n15225), .A2(n14864), .B1(n15226), .C1(n15227), .Y(
        n15224) );
  a21oi_1 U14200 ( .A1(n15009), .A2(n15228), .B1(n14850), .Y(n15227) );
  inv_1 U14201 ( .A(n15131), .Y(n15225) );
  inv_1 U14202 ( .A(n15229), .Y(n15223) );
  or3_1 U14203 ( .A(n15115), .B(n15230), .C(n15231), .X(n14932) );
  o221ai_1 U14204 ( .A1(n15086), .A2(n14848), .B1(n14880), .B2(n15076), .C1(
        n15037), .Y(n15231) );
  inv_1 U14205 ( .A(n15232), .Y(n15230) );
  o22ai_1 U14206 ( .A1(n15233), .A2(n14848), .B1(n15234), .B2(n14997), .Y(
        n15115) );
  nand2_1 U14207 ( .A(n14941), .B(n15124), .Y(n15221) );
  inv_1 U14208 ( .A(n15235), .Y(n15124) );
  o21ai_0 U14209 ( .A1(n15236), .A2(n14897), .B1(n15237), .Y(n15235) );
  a21oi_1 U14210 ( .A1(n14864), .A2(n15238), .B1(n15239), .Y(n14941) );
  nor4_1 U14211 ( .A(n15119), .B(n15079), .C(n15138), .D(n15190), .Y(n15191)
         );
  o221ai_1 U14212 ( .A1(n15240), .A2(n14895), .B1(n14997), .B2(n15241), .C1(
        n15129), .Y(n15190) );
  nand3_1 U14213 ( .A(n15242), .B(n15200), .C(n14922), .Y(n15129) );
  and3_1 U14214 ( .A(n15010), .B(n15032), .C(n14878), .X(n15240) );
  nand2_1 U14215 ( .A(n12461), .B(n15243), .Y(n14878) );
  o22ai_1 U14216 ( .A1(n14895), .A2(n15034), .B1(n15244), .B2(n14942), .Y(
        n15138) );
  inv_1 U14217 ( .A(n15182), .Y(n15244) );
  or3_1 U14218 ( .A(n15245), .B(n14951), .C(n15246), .X(n15079) );
  inv_1 U14219 ( .A(n15247), .Y(n15246) );
  a211oi_1 U14220 ( .A1(n15248), .A2(n14965), .B1(n15097), .C1(n15249), .Y(
        n15247) );
  and3_1 U14221 ( .A(n14946), .B(n15250), .C(n15251), .X(n15097) );
  nand2_1 U14222 ( .A(n15252), .B(n15253), .Y(n14951) );
  o21ai_0 U14223 ( .A1(n15254), .A2(n15255), .B1(n14986), .Y(n15253) );
  inv_1 U14224 ( .A(n15122), .Y(n15255) );
  nor4_1 U14225 ( .A(n15256), .B(n15180), .C(n15257), .D(n15258), .Y(n15254)
         );
  o32ai_1 U14226 ( .A1(n15076), .A2(n14960), .A3(n15259), .B1(n15260), .B2(
        n12466), .Y(n15119) );
  nor2_1 U14227 ( .A(n14856), .B(n15261), .Y(n15260) );
  or4_1 U14228 ( .A(n15039), .B(n15189), .C(n15262), .D(n15263), .X(n10366) );
  nand4_1 U14229 ( .A(n12458), .B(n15264), .C(n15265), .D(n15266), .Y(n15263)
         );
  a222oi_1 U14230 ( .A1(n15016), .A2(n14946), .B1(n15267), .B2(n14964), .C1(
        n14908), .C2(n14887), .Y(n15266) );
  nand2_1 U14231 ( .A(n15268), .B(n15004), .Y(n14887) );
  inv_1 U14232 ( .A(n15174), .Y(n15004) );
  nor2_1 U14233 ( .A(n15202), .B(n14962), .Y(n15174) );
  nand4_1 U14234 ( .A(n15023), .B(n15269), .C(n15117), .D(n15270), .Y(n15267)
         );
  a21oi_1 U14235 ( .A1(n12461), .A2(n14873), .B1(n14888), .Y(n15270) );
  nand2_1 U14236 ( .A(n14998), .B(n15050), .Y(n14888) );
  nand3_1 U14237 ( .A(n14872), .B(n12462), .C(n15271), .Y(n15050) );
  nand4_1 U14238 ( .A(n15205), .B(n15272), .C(n14919), .D(n15214), .Y(n15117)
         );
  inv_1 U14239 ( .A(n15179), .Y(n15016) );
  o21ai_0 U14240 ( .A1(n15273), .A2(n14892), .B1(n14922), .Y(n15265) );
  nand2_1 U14241 ( .A(n15274), .B(n14943), .Y(n14892) );
  nand3_1 U14242 ( .A(n15025), .B(n14901), .C(n15275), .Y(n15262) );
  inv_1 U14243 ( .A(n14929), .Y(n15275) );
  o22ai_1 U14244 ( .A1(n12466), .A2(n15276), .B1(n14859), .B2(n15036), .Y(
        n14929) );
  nor4_1 U14245 ( .A(n15165), .B(n15222), .C(n15277), .D(n15278), .Y(n14901)
         );
  inv_1 U14246 ( .A(n15279), .Y(n15278) );
  a211oi_1 U14247 ( .A1(n15006), .A2(n14908), .B1(n15280), .C1(n15022), .Y(
        n15279) );
  o211ai_1 U14248 ( .A1(n12466), .A2(n15206), .B1(n15281), .C1(n15282), .Y(
        n15022) );
  a211oi_1 U14249 ( .A1(n15283), .A2(n12460), .B1(n15284), .C1(n15144), .Y(
        n15282) );
  inv_1 U14250 ( .A(n12459), .Y(n15144) );
  inv_1 U14251 ( .A(n15219), .Y(n15281) );
  o21ai_0 U14252 ( .A1(n12466), .A2(n14970), .B1(n15285), .Y(n15219) );
  o21ai_0 U14253 ( .A1(n12466), .A2(n15049), .B1(n15166), .Y(n15280) );
  nand2_1 U14254 ( .A(n15286), .B(n15102), .Y(n15166) );
  inv_1 U14255 ( .A(n14897), .Y(n14908) );
  inv_1 U14256 ( .A(n15241), .Y(n15006) );
  or3_1 U14257 ( .A(n15132), .B(n15287), .C(n15065), .X(n15222) );
  nor4_1 U14258 ( .A(n15288), .B(n15258), .C(n15257), .D(n14997), .Y(n15065)
         );
  inv_1 U14259 ( .A(n15024), .Y(n15287) );
  nand4_1 U14260 ( .A(n15289), .B(n15250), .C(n15290), .D(n14965), .Y(n15024)
         );
  nor2_1 U14261 ( .A(n15291), .B(n12466), .Y(n15132) );
  or4_1 U14262 ( .A(n15098), .B(n15249), .C(n14959), .D(n15239), .X(n15165) );
  nor3_1 U14263 ( .A(n15076), .B(n14984), .C(n15202), .Y(n15239) );
  a211oi_1 U14264 ( .A1(n15292), .A2(n15067), .B1(n14897), .C1(n15068), .Y(
        n15098) );
  a221oi_1 U14265 ( .A1(n15293), .A2(n14965), .B1(n14988), .B2(n12460), .C1(
        n15294), .Y(n15025) );
  nand2_1 U14266 ( .A(n15295), .B(n15149), .Y(n15293) );
  o221ai_1 U14267 ( .A1(n12466), .A2(n14917), .B1(n15076), .B2(n15296), .C1(
        n15297), .Y(n15189) );
  inv_1 U14268 ( .A(n15298), .Y(n15297) );
  o221ai_1 U14269 ( .A1(n15228), .A2(n14850), .B1(n15299), .B2(n14859), .C1(
        n15037), .Y(n15298) );
  and3_1 U14270 ( .A(n14870), .B(n14881), .C(n15122), .X(n15299) );
  nand3_1 U14271 ( .A(n15300), .B(n15158), .C(n15161), .Y(n15122) );
  nand2_1 U14272 ( .A(n15301), .B(n15302), .Y(n15228) );
  o32ai_1 U14273 ( .A1(n15303), .A2(n15304), .A3(n15305), .B1(n15306), .B2(
        n15307), .Y(n15302) );
  nand2_1 U14274 ( .A(n15215), .B(n15308), .Y(n14917) );
  nand3_1 U14275 ( .A(n15232), .B(n15309), .C(n15310), .Y(n15039) );
  nor3_1 U14276 ( .A(n15127), .B(n15096), .C(n15226), .Y(n15310) );
  and4_1 U14277 ( .A(n23873), .B(n15311), .C(n15243), .D(n15312), .X(n15226)
         );
  nor3_1 U14278 ( .A(n15303), .B(n14889), .C(n14850), .Y(n15312) );
  inv_1 U14279 ( .A(n15167), .Y(n15096) );
  nand4_1 U14280 ( .A(n14986), .B(n15313), .C(n15314), .D(n15315), .Y(n15167)
         );
  o32ai_1 U14281 ( .A1(n14982), .A2(n15256), .A3(n15180), .B1(n15316), .B2(
        n15288), .Y(n15315) );
  o21ai_0 U14282 ( .A1(n15238), .A2(n15182), .B1(n14864), .Y(n15309) );
  nand2_1 U14283 ( .A(n15062), .B(n14894), .Y(n15182) );
  nand3_1 U14284 ( .A(n15213), .B(n15301), .C(n15317), .Y(n15062) );
  a21oi_1 U14285 ( .A1(n14986), .A2(n15318), .B1(n15128), .Y(n15232) );
  and4_1 U14286 ( .A(n15158), .B(n23873), .C(n15319), .D(n15320), .X(n15128)
         );
  nor2_1 U14287 ( .A(n14895), .B(n15307), .Y(n15320) );
  and2_0 U14288 ( .A(n15321), .B(n10614), .X(n15318) );
  nand3_1 U14289 ( .A(n15322), .B(n15323), .C(n15324), .Y(n10365) );
  nor4_1 U14290 ( .A(n15325), .B(n15326), .C(n14959), .D(n15294), .Y(n15324)
         );
  and4_1 U14291 ( .A(n15319), .B(n15327), .C(n15328), .D(n15329), .X(n15294)
         );
  nor3_1 U14292 ( .A(n14895), .B(n15330), .C(n15292), .Y(n15329) );
  nor2_1 U14293 ( .A(n15121), .B(n15076), .Y(n14959) );
  a21oi_1 U14294 ( .A1(n15331), .A2(n15157), .B1(n14942), .Y(n15326) );
  nand4_1 U14295 ( .A(n15237), .B(n15332), .C(n15333), .D(n15285), .Y(n15325)
         );
  nand4_1 U14296 ( .A(n14855), .B(n23873), .C(n15334), .D(n15335), .Y(n15285)
         );
  nor2_1 U14297 ( .A(n15303), .B(n14848), .Y(n15335) );
  inv_1 U14298 ( .A(n14846), .Y(n15332) );
  nor3_1 U14299 ( .A(n15202), .B(n15203), .C(n14942), .Y(n14846) );
  or2_0 U14300 ( .A(n15013), .B(n14942), .X(n15237) );
  nor3_1 U14301 ( .A(n15336), .B(n15229), .C(n14930), .Y(n15323) );
  or3_1 U14302 ( .A(n14945), .B(n15337), .C(n15338), .X(n14930) );
  o211ai_1 U14303 ( .A1(n15009), .A2(n14850), .B1(n15264), .C1(n15339), .Y(
        n15338) );
  o22ai_1 U14304 ( .A1(n12463), .A2(n14848), .B1(n14897), .B2(n15150), .Y(
        n14945) );
  o22ai_1 U14305 ( .A1(n14850), .A2(n14918), .B1(n15076), .B2(n15077), .Y(
        n15229) );
  o22ai_1 U14306 ( .A1(n14859), .A2(n15340), .B1(n15236), .B2(n14997), .Y(
        n15336) );
  and2_0 U14307 ( .A(n15172), .B(n14881), .X(n15236) );
  nor4_1 U14308 ( .A(n15341), .B(n15342), .C(n14853), .D(n15343), .Y(n15340)
         );
  inv_1 U14309 ( .A(n15051), .Y(n14853) );
  nand3_1 U14310 ( .A(n15344), .B(n15216), .C(n14998), .Y(n15342) );
  nand3_1 U14311 ( .A(n14909), .B(n15304), .C(n14852), .Y(n15216) );
  nand4_1 U14312 ( .A(n15345), .B(n14977), .C(n15346), .D(n15296), .Y(n15341)
         );
  and4_1 U14313 ( .A(n15052), .B(n15071), .C(n15347), .D(n14880), .X(n14977)
         );
  inv_1 U14314 ( .A(n15348), .Y(n15345) );
  nor3_1 U14315 ( .A(n15349), .B(n15139), .C(n15176), .Y(n15322) );
  o22ai_1 U14316 ( .A1(n14897), .A2(n15036), .B1(n14848), .B2(n15049), .Y(
        n15176) );
  nand3_1 U14317 ( .A(n15317), .B(n15242), .C(n15205), .Y(n15049) );
  o22ai_1 U14318 ( .A1(n14848), .A2(n15179), .B1(n14897), .B2(n15241), .Y(
        n15139) );
  nand3_1 U14319 ( .A(n15350), .B(n15351), .C(n15352), .Y(n10364) );
  nor4_1 U14320 ( .A(n15353), .B(n15354), .C(n15355), .D(n15356), .Y(n15352)
         );
  a21oi_1 U14321 ( .A1(n15234), .A2(n15268), .B1(n14897), .Y(n15356) );
  and4_1 U14322 ( .A(n15150), .B(n14996), .C(n15075), .D(n15057), .X(n15268)
         );
  nand2_1 U14323 ( .A(n15215), .B(n14851), .Y(n14996) );
  and3_1 U14324 ( .A(n15243), .B(n15357), .C(n15358), .X(n15215) );
  nand3_1 U14325 ( .A(n15359), .B(n14920), .C(n15358), .Y(n15150) );
  inv_1 U14326 ( .A(n15059), .Y(n15234) );
  o21ai_0 U14327 ( .A1(n14973), .A2(n14962), .B1(n15360), .Y(n15059) );
  a21oi_1 U14328 ( .A1(n15034), .A2(n15269), .B1(n14942), .Y(n15355) );
  nand3_1 U14329 ( .A(n15205), .B(n15204), .C(n14874), .Y(n15269) );
  inv_1 U14330 ( .A(n14981), .Y(n14874) );
  o22ai_1 U14331 ( .A1(n14859), .A2(n15361), .B1(n14850), .B2(n14880), .Y(
        n15354) );
  nand4_1 U14332 ( .A(n23892), .B(n15362), .C(n15363), .D(n15364), .Y(n14880)
         );
  nor2_1 U14333 ( .A(n15259), .B(n15365), .Y(n15364) );
  nor4_1 U14334 ( .A(n15366), .B(n15367), .C(n15348), .D(n15368), .Y(n15361)
         );
  o21ai_0 U14335 ( .A1(n15068), .A2(n14981), .B1(n15369), .Y(n15368) );
  inv_1 U14336 ( .A(n15110), .Y(n15369) );
  nand3_1 U14337 ( .A(n14870), .B(n15032), .C(n15155), .Y(n15110) );
  inv_1 U14338 ( .A(n14923), .Y(n15155) );
  nand2_1 U14339 ( .A(n14943), .B(n15023), .Y(n14923) );
  inv_1 U14340 ( .A(n14863), .Y(n15023) );
  nor4_1 U14341 ( .A(n15303), .B(n14889), .C(n14968), .D(n15370), .Y(n14863)
         );
  nand2_1 U14342 ( .A(n15251), .B(n15242), .Y(n14870) );
  inv_1 U14343 ( .A(n14889), .Y(n15242) );
  nand2_1 U14344 ( .A(n15371), .B(n15372), .Y(n14981) );
  nand3_1 U14345 ( .A(n15030), .B(n15087), .C(n15108), .Y(n15348) );
  inv_1 U14346 ( .A(n15248), .Y(n15030) );
  nor2_1 U14347 ( .A(n15068), .B(n15292), .Y(n15248) );
  nand3_1 U14348 ( .A(n15241), .B(n15077), .C(n15291), .Y(n15367) );
  nand4_1 U14349 ( .A(n15373), .B(n15374), .C(n15375), .D(n15376), .Y(n15241)
         );
  nor4_1 U14350 ( .A(n23922), .B(n23892), .C(n23871), .D(n14873), .Y(n15376)
         );
  nand4_1 U14351 ( .A(n15347), .B(n15152), .C(n15131), .D(n15377), .Y(n15366)
         );
  and3_1 U14352 ( .A(n14881), .B(n15157), .C(n15121), .X(n15377) );
  nand3_1 U14353 ( .A(n15158), .B(n15378), .C(n15379), .Y(n15121) );
  nand2_1 U14354 ( .A(n14921), .B(n15378), .Y(n14881) );
  nand2_1 U14355 ( .A(n15250), .B(n15200), .Y(n15131) );
  inv_1 U14356 ( .A(n14856), .Y(n15347) );
  nor2_1 U14357 ( .A(n15151), .B(n10614), .Y(n14856) );
  nand4_1 U14358 ( .A(n15380), .B(n15037), .C(n15199), .D(n15136), .Y(n15353)
         );
  nand4_1 U14359 ( .A(n15272), .B(n15271), .C(n14986), .D(n15301), .Y(n15136)
         );
  nand4_1 U14360 ( .A(n14922), .B(n15204), .C(n15381), .D(n15301), .Y(n15037)
         );
  o21ai_0 U14361 ( .A1(n15261), .A2(n15382), .B1(n14946), .Y(n15380) );
  inv_1 U14362 ( .A(n14970), .Y(n15382) );
  nand3_1 U14363 ( .A(n15378), .B(n15383), .C(n15379), .Y(n14970) );
  nor2_1 U14364 ( .A(n14857), .B(n15008), .Y(n15261) );
  nand4_1 U14365 ( .A(n15185), .B(n15327), .C(n23893), .D(n10614), .Y(n14857)
         );
  nor3_1 U14366 ( .A(n15384), .B(n15277), .C(n15385), .Y(n15351) );
  inv_1 U14367 ( .A(n14840), .Y(n15385) );
  nor4_1 U14368 ( .A(n15074), .B(n15066), .C(n15386), .D(n15387), .Y(n14840)
         );
  o221ai_1 U14369 ( .A1(n15011), .A2(n12466), .B1(n15172), .B2(n14997), .C1(
        n15175), .Y(n15387) );
  nor3_1 U14370 ( .A(n15388), .B(n14955), .C(n15127), .Y(n15175) );
  inv_1 U14371 ( .A(n15339), .Y(n15127) );
  nand4_1 U14372 ( .A(n15389), .B(n15362), .C(n15390), .D(n15391), .Y(n15339)
         );
  nor3_1 U14373 ( .A(n14850), .B(n15258), .C(n15292), .Y(n15391) );
  and3_1 U14374 ( .A(n15321), .B(n12462), .C(n14986), .X(n14955) );
  inv_1 U14375 ( .A(n15264), .Y(n15388) );
  nand3_1 U14376 ( .A(n12461), .B(n12462), .C(n14986), .Y(n15264) );
  nand2_1 U14377 ( .A(n12461), .B(n15300), .Y(n15172) );
  inv_1 U14378 ( .A(n15130), .Y(n15011) );
  nor2_1 U14379 ( .A(n15151), .B(n23837), .Y(n15130) );
  o21ai_0 U14380 ( .A1(n15013), .A2(n14895), .B1(n15252), .Y(n15386) );
  nand2_1 U14381 ( .A(n14851), .B(n15392), .Y(n15013) );
  nor3_1 U14382 ( .A(n14942), .B(n15007), .C(n14889), .Y(n15066) );
  nand2_1 U14383 ( .A(n15393), .B(n15394), .Y(n14889) );
  nor2_1 U14384 ( .A(n15163), .B(n12466), .Y(n15074) );
  o221ai_1 U14385 ( .A1(n12466), .A2(n15052), .B1(n15162), .B2(n14848), .C1(
        n15073), .Y(n15277) );
  nand4_1 U14386 ( .A(n15161), .B(n14946), .C(n14851), .D(n15378), .Y(n15073)
         );
  and4_1 U14387 ( .A(n15233), .B(n15395), .C(n15086), .D(n12463), .X(n15162)
         );
  nand3_1 U14388 ( .A(n15334), .B(n15250), .C(n15396), .Y(n12463) );
  nor3_1 U14389 ( .A(n15258), .B(n23873), .C(n15256), .Y(n15396) );
  nand3_1 U14390 ( .A(n14851), .B(n12462), .C(n15397), .Y(n15086) );
  nand2_1 U14391 ( .A(n15251), .B(n15250), .Y(n15395) );
  and4_1 U14392 ( .A(n15390), .B(n15398), .C(n15375), .D(n15399), .X(n15251)
         );
  nor3_1 U14393 ( .A(n23873), .B(n23922), .C(n23892), .Y(n15399) );
  a21oi_1 U14394 ( .A1(n15378), .A2(n12461), .B1(n15400), .Y(n15233) );
  and4_1 U14395 ( .A(n15308), .B(n15204), .C(n15390), .D(n15362), .X(n15400)
         );
  inv_1 U14396 ( .A(n14969), .Y(n12461) );
  nand2_1 U14397 ( .A(n15308), .B(n15397), .Y(n14969) );
  and3_1 U14398 ( .A(n23873), .B(n15311), .C(n15204), .X(n15397) );
  nand3_1 U14399 ( .A(n15401), .B(n15314), .C(n15317), .Y(n15052) );
  inv_1 U14400 ( .A(n15102), .Y(n12466) );
  o22ai_1 U14401 ( .A1(n14895), .A2(n15091), .B1(n15076), .B2(n15009), .Y(
        n15384) );
  nor3_1 U14402 ( .A(n15188), .B(n15080), .C(n15137), .Y(n15350) );
  or3_1 U14403 ( .A(n15249), .B(n15284), .C(n15402), .X(n15137) );
  a21oi_1 U14404 ( .A1(n15295), .A2(n15036), .B1(n14997), .Y(n15402) );
  nand4_1 U14405 ( .A(n15204), .B(n15213), .C(n12462), .D(n15314), .Y(n15036)
         );
  inv_1 U14406 ( .A(n15333), .Y(n15284) );
  nand4_1 U14407 ( .A(n15205), .B(n15272), .C(n15383), .D(n14965), .Y(n15333)
         );
  and3_1 U14408 ( .A(n15272), .B(n15213), .C(n15403), .X(n15249) );
  nor3_1 U14409 ( .A(n14968), .B(n15370), .C(n14997), .Y(n15403) );
  o221ai_1 U14410 ( .A1(n15404), .A2(n14942), .B1(n15076), .B2(n14998), .C1(
        n15405), .Y(n15080) );
  a21oi_1 U14411 ( .A1(n14986), .A2(n15406), .B1(n15407), .Y(n15405) );
  inv_1 U14412 ( .A(n15408), .Y(n15407) );
  o211ai_1 U14413 ( .A1(n14984), .A2(n15202), .B1(n15296), .C1(n15135), .Y(
        n15406) );
  nand3_1 U14414 ( .A(n15308), .B(n15301), .C(n15409), .Y(n15135) );
  inv_1 U14415 ( .A(n15303), .Y(n15409) );
  nand2_1 U14416 ( .A(n15290), .B(n15410), .Y(n15303) );
  inv_1 U14417 ( .A(n15256), .Y(n15290) );
  nand4_1 U14418 ( .A(n15358), .B(n15271), .C(n12462), .D(n15357), .Y(n15296)
         );
  inv_1 U14419 ( .A(n15411), .Y(n15358) );
  nand3_1 U14420 ( .A(n15272), .B(n15373), .C(n15205), .Y(n14998) );
  inv_1 U14421 ( .A(n14914), .Y(n15404) );
  nand2_1 U14422 ( .A(n14871), .B(n14894), .Y(n14914) );
  nand4_1 U14423 ( .A(n15412), .B(n15413), .C(n15393), .D(n15371), .Y(n14894)
         );
  o221ai_1 U14424 ( .A1(n15414), .A2(n14848), .B1(n14884), .B2(n15076), .C1(
        n15100), .Y(n15188) );
  inv_1 U14425 ( .A(n14987), .Y(n14884) );
  o21ai_0 U14426 ( .A1(n15007), .A2(n15180), .B1(n15220), .Y(n14987) );
  and2_0 U14427 ( .A(n15206), .B(n15058), .X(n15414) );
  nand4_1 U14428 ( .A(n15415), .B(n15416), .C(n15417), .D(n15418), .Y(n10363)
         );
  nor4_1 U14429 ( .A(n14907), .B(n15419), .C(n15420), .D(n15421), .Y(n15418)
         );
  a21oi_1 U14430 ( .A1(n15091), .A2(n15163), .B1(n14859), .Y(n15421) );
  nand4_1 U14431 ( .A(n15317), .B(n14855), .C(n15300), .D(n15314), .Y(n15163)
         );
  nand4_1 U14432 ( .A(n12462), .B(n15314), .C(n15250), .D(n15422), .Y(n15091)
         );
  nor2_1 U14433 ( .A(n15330), .B(n15411), .Y(n15422) );
  nand2_1 U14434 ( .A(n15328), .B(n23892), .Y(n15411) );
  and2_0 U14435 ( .A(n15371), .B(n14919), .X(n15250) );
  inv_1 U14436 ( .A(n12458), .Y(n15420) );
  nand2_1 U14437 ( .A(n14964), .B(n15423), .Y(n12458) );
  nand4_1 U14438 ( .A(n15424), .B(n14858), .C(n15346), .D(n15425), .Y(n15423)
         );
  inv_1 U14439 ( .A(n15426), .Y(n15425) );
  o211ai_1 U14440 ( .A1(n15114), .A2(n14960), .B1(n15157), .C1(n15151), .Y(
        n15426) );
  nand4_1 U14441 ( .A(n15185), .B(n15158), .C(n15314), .D(n23892), .Y(n15151)
         );
  nand4_1 U14442 ( .A(n15378), .B(n15383), .C(n14876), .D(n15311), .Y(n15157)
         );
  nand2_1 U14443 ( .A(n14909), .B(n15427), .Y(n15114) );
  and4_1 U14444 ( .A(n14879), .B(n15152), .C(n15012), .D(n15428), .X(n15346)
         );
  nor3_1 U14445 ( .A(n15061), .B(n15089), .C(n15429), .Y(n15428) );
  nor4_1 U14446 ( .A(n15311), .B(n15430), .C(n15113), .D(n15008), .Y(n15429)
         );
  nand2_1 U14447 ( .A(n23872), .B(n15394), .Y(n15008) );
  inv_1 U14448 ( .A(n15220), .Y(n15089) );
  nand4_1 U14449 ( .A(n15301), .B(n15383), .C(n15431), .D(n15184), .Y(n15220)
         );
  inv_1 U14450 ( .A(n15203), .Y(n15383) );
  and2_0 U14451 ( .A(n15390), .B(n23873), .X(n15301) );
  nand4_1 U14452 ( .A(n15432), .B(n14896), .C(n15010), .D(n15034), .Y(n15061)
         );
  nand3_1 U14453 ( .A(n14877), .B(n14876), .C(n15319), .Y(n15034) );
  nand4_1 U14454 ( .A(n15401), .B(n15363), .C(n15327), .D(n15311), .Y(n15010)
         );
  and3_1 U14455 ( .A(n15371), .B(n15300), .C(n15393), .X(n15401) );
  nand4_1 U14456 ( .A(n15374), .B(n15185), .C(n15158), .D(n15184), .Y(n14896)
         );
  nand4_1 U14457 ( .A(n14855), .B(n14875), .C(n15185), .D(n23873), .Y(n15432)
         );
  nand3_1 U14458 ( .A(n15200), .B(n15433), .C(n14919), .Y(n15012) );
  inv_1 U14459 ( .A(n15007), .Y(n15200) );
  nand3_1 U14460 ( .A(n15185), .B(n15327), .C(n14875), .Y(n15007) );
  inv_1 U14461 ( .A(n15187), .Y(n14875) );
  nand3_1 U14462 ( .A(n14852), .B(n23894), .C(n15359), .Y(n15152) );
  inv_1 U14463 ( .A(n14960), .Y(n14852) );
  nand2_1 U14464 ( .A(n15390), .B(n14876), .Y(n14960) );
  nor2_1 U14465 ( .A(n15187), .B(n14873), .Y(n15390) );
  nand3_1 U14466 ( .A(n14909), .B(n24036), .C(n15392), .Y(n14879) );
  inv_1 U14467 ( .A(n14973), .Y(n15392) );
  nand3_1 U14468 ( .A(n15185), .B(n23892), .C(n15374), .Y(n14973) );
  inv_1 U14469 ( .A(n15113), .Y(n15185) );
  nand2_1 U14470 ( .A(n15363), .B(n24037), .Y(n15113) );
  and2_0 U14471 ( .A(n15071), .B(n15087), .X(n14858) );
  nand4_1 U14472 ( .A(n15213), .B(n15300), .C(n14876), .D(n15311), .Y(n15087)
         );
  and2_0 U14473 ( .A(n15327), .B(n15431), .X(n14876) );
  nand4_1 U14474 ( .A(n15431), .B(n23873), .C(n15158), .D(n15434), .Y(n15071)
         );
  and3_1 U14475 ( .A(n12462), .B(n15184), .C(n23893), .X(n15434) );
  inv_1 U14476 ( .A(n14984), .Y(n15158) );
  nand2_1 U14477 ( .A(n15214), .B(n14909), .Y(n14984) );
  nor3_1 U14478 ( .A(n15256), .B(n10774), .C(n15435), .Y(n15431) );
  nand2_1 U14479 ( .A(n23836), .B(n15398), .Y(n15256) );
  inv_1 U14480 ( .A(n15159), .Y(n15424) );
  nand2_1 U14481 ( .A(n15009), .B(n15436), .Y(n15159) );
  nand4_1 U14482 ( .A(n14851), .B(n15374), .C(n15363), .D(n23892), .Y(n15436)
         );
  inv_1 U14483 ( .A(n15112), .Y(n15374) );
  nand3_1 U14484 ( .A(n10614), .B(n15362), .C(n23893), .Y(n15112) );
  nand4_1 U14485 ( .A(n15381), .B(n15437), .C(n15363), .D(n23892), .Y(n15009)
         );
  and3_1 U14486 ( .A(n23838), .B(n23922), .C(n15389), .X(n15363) );
  inv_1 U14487 ( .A(n15199), .Y(n15419) );
  nand2_1 U14488 ( .A(n15343), .B(n14946), .Y(n15199) );
  inv_1 U14489 ( .A(n15276), .Y(n15343) );
  nand3_1 U14490 ( .A(n15213), .B(n12462), .C(n15161), .Y(n15276) );
  nor3_1 U14491 ( .A(n14848), .B(n14982), .C(n15085), .Y(n14907) );
  a222oi_1 U14492 ( .A1(n15238), .A2(n14922), .B1(n15102), .B2(n14985), .C1(
        n14986), .C2(n14988), .Y(n15417) );
  nand2_1 U14493 ( .A(n15051), .B(n15077), .Y(n14988) );
  nand3_1 U14494 ( .A(n15381), .B(n15300), .C(n15379), .Y(n15077) );
  inv_1 U14495 ( .A(n14962), .Y(n15381) );
  nand4_1 U14496 ( .A(n14925), .B(n15313), .C(n15378), .D(n15357), .Y(n15051)
         );
  inv_1 U14497 ( .A(n14968), .Y(n15378) );
  nand2_1 U14498 ( .A(n23837), .B(n24037), .Y(n14968) );
  nand2_1 U14499 ( .A(n15179), .B(n15058), .Y(n14985) );
  nand4_1 U14500 ( .A(n15317), .B(n15334), .C(n14877), .D(n23873), .Y(n15058)
         );
  nor2_1 U14501 ( .A(n15330), .B(n15438), .Y(n15317) );
  nand2_1 U14502 ( .A(n14921), .B(n15300), .Y(n15179) );
  inv_1 U14503 ( .A(n15316), .Y(n15300) );
  nand2_1 U14504 ( .A(n23837), .B(n14873), .Y(n15316) );
  inv_1 U14505 ( .A(n15085), .Y(n14921) );
  nand3_1 U14506 ( .A(n14877), .B(n15314), .C(n15204), .Y(n15085) );
  nor2_1 U14507 ( .A(n15439), .B(n14859), .Y(n15102) );
  inv_1 U14508 ( .A(n14871), .Y(n15238) );
  nand3_1 U14509 ( .A(n14925), .B(n12462), .C(n15161), .Y(n14871) );
  and4_1 U14510 ( .A(n15413), .B(n15328), .C(n15327), .D(n15311), .X(n15161)
         );
  inv_1 U14511 ( .A(n15440), .Y(n14925) );
  a211oi_1 U14512 ( .A1(n15441), .A2(n14946), .B1(n14940), .C1(n15337), .Y(
        n15416) );
  o21ai_0 U14513 ( .A1(n14848), .A2(n15206), .B1(n15408), .Y(n15337) );
  nand2_1 U14514 ( .A(n15283), .B(n14986), .Y(n15408) );
  inv_1 U14515 ( .A(n14850), .Y(n14986) );
  nand2_1 U14516 ( .A(n15442), .B(n14964), .Y(n14850) );
  and4_1 U14517 ( .A(n15313), .B(n15243), .C(n14877), .D(n15357), .X(n15283)
         );
  inv_1 U14518 ( .A(n15217), .Y(n14877) );
  nand2_1 U14519 ( .A(n15359), .B(n15394), .Y(n15217) );
  nand3_1 U14520 ( .A(n15359), .B(n14920), .C(n15313), .Y(n15206) );
  o221ai_1 U14521 ( .A1(n14942), .A2(n15032), .B1(n15076), .B2(n14918), .C1(
        n15100), .Y(n14940) );
  nand2_1 U14522 ( .A(n14864), .B(n15443), .Y(n15100) );
  o21ai_0 U14523 ( .A1(n15203), .A2(n15202), .B1(n15274), .Y(n15443) );
  nor2_1 U14524 ( .A(n15090), .B(n15017), .Y(n15274) );
  and3_1 U14525 ( .A(n15308), .B(n15389), .C(n15412), .X(n15017) );
  and3_1 U14526 ( .A(n12462), .B(n15314), .C(n15313), .X(n15412) );
  nor2_1 U14527 ( .A(n15305), .B(n14961), .Y(n15308) );
  inv_1 U14528 ( .A(n15214), .Y(n14961) );
  inv_1 U14529 ( .A(n15331), .Y(n15090) );
  nand4_1 U14530 ( .A(n15271), .B(n15204), .C(n15319), .D(n23873), .Y(n15331)
         );
  inv_1 U14531 ( .A(n15306), .Y(n15271) );
  nand4_1 U14532 ( .A(n15328), .B(n15243), .C(n15357), .D(n15184), .Y(n15202)
         );
  nand2_1 U14533 ( .A(n15394), .B(n14909), .Y(n15203) );
  inv_1 U14534 ( .A(n15021), .Y(n14918) );
  nor2_1 U14535 ( .A(n15306), .B(n15068), .Y(n15021) );
  nand2_1 U14536 ( .A(n14919), .B(n15444), .Y(n15306) );
  inv_1 U14537 ( .A(n15273), .Y(n15032) );
  nor2_1 U14538 ( .A(n14891), .B(n15258), .Y(n15273) );
  nand4_1 U14539 ( .A(n15334), .B(n15213), .C(n15389), .D(n15362), .Y(n14891)
         );
  inv_1 U14540 ( .A(n15365), .Y(n15334) );
  inv_1 U14541 ( .A(n14848), .Y(n14946) );
  inv_1 U14542 ( .A(n15291), .Y(n15441) );
  nand3_1 U14543 ( .A(n15437), .B(n14855), .C(n15272), .Y(n15291) );
  inv_1 U14544 ( .A(n15307), .Y(n15272) );
  nand3_1 U14545 ( .A(n15328), .B(n15184), .C(n15413), .Y(n15307) );
  inv_1 U14546 ( .A(n15330), .Y(n15413) );
  nand2_1 U14547 ( .A(n23871), .B(n15445), .Y(n15330) );
  nor2_1 U14548 ( .A(n15435), .B(n23922), .Y(n15328) );
  inv_1 U14549 ( .A(n15180), .Y(n14855) );
  nand2_1 U14550 ( .A(n14919), .B(n15394), .Y(n15180) );
  inv_1 U14551 ( .A(n15427), .Y(n15394) );
  nand2_1 U14552 ( .A(n23894), .B(n15433), .Y(n15427) );
  inv_1 U14553 ( .A(n15257), .Y(n15437) );
  nand2_1 U14554 ( .A(n15243), .B(n15314), .Y(n15257) );
  inv_1 U14555 ( .A(n15370), .Y(n15314) );
  nor3_1 U14556 ( .A(n15349), .B(n15245), .C(n15177), .Y(n15415) );
  o21ai_0 U14557 ( .A1(n15076), .A2(n15108), .B1(n15038), .Y(n15177) );
  nand3_1 U14558 ( .A(n14922), .B(n15289), .C(n15446), .Y(n15038) );
  inv_1 U14559 ( .A(n15288), .Y(n15446) );
  nand3_1 U14560 ( .A(n15214), .B(n15389), .C(n14919), .Y(n15288) );
  inv_1 U14561 ( .A(n14895), .Y(n14922) );
  nand2_1 U14562 ( .A(n15447), .B(n14964), .Y(n14895) );
  nand2_1 U14563 ( .A(n15321), .B(n15243), .Y(n15108) );
  nor2_1 U14564 ( .A(n15440), .B(n14983), .Y(n15321) );
  inv_1 U14565 ( .A(n12460), .Y(n15076) );
  nor2_1 U14566 ( .A(n15442), .B(n14859), .Y(n12460) );
  nor2_1 U14567 ( .A(n15448), .B(inData[23]), .Y(n15442) );
  o22ai_1 U14568 ( .A1(n14897), .A2(n15295), .B1(n15344), .B2(n14848), .Y(
        n15245) );
  nand2_1 U14569 ( .A(n15439), .B(n14964), .Y(n14848) );
  nor2_1 U14570 ( .A(n15449), .B(n15448), .Y(n15439) );
  inv_1 U14571 ( .A(n15286), .Y(n15344) );
  nor2_1 U14572 ( .A(n15068), .B(n15440), .Y(n15286) );
  nand2_1 U14573 ( .A(n15371), .B(n14909), .Y(n15440) );
  nand2_1 U14574 ( .A(n15379), .B(n15243), .Y(n15068) );
  and2_0 U14575 ( .A(n15410), .B(n15357), .X(n15379) );
  nand3_1 U14576 ( .A(n15213), .B(n15243), .C(n14872), .Y(n15295) );
  inv_1 U14577 ( .A(n14983), .Y(n14872) );
  nand3_1 U14578 ( .A(n23893), .B(n15362), .C(n15204), .Y(n14983) );
  and2_0 U14579 ( .A(n15389), .B(n15410), .X(n15204) );
  inv_1 U14580 ( .A(n15067), .Y(n15213) );
  nand2_1 U14581 ( .A(n15371), .B(n15359), .Y(n15067) );
  nor2_1 U14582 ( .A(n23894), .B(n24036), .Y(n15371) );
  nand4_1 U14583 ( .A(n15450), .B(n15451), .C(n15252), .D(n12459), .Y(n15349)
         );
  nand2_1 U14584 ( .A(n14965), .B(n15452), .Y(n12459) );
  or2_0 U14585 ( .A(n15149), .B(n14897), .X(n15252) );
  nand2_1 U14586 ( .A(n15453), .B(n14964), .Y(n14897) );
  nand3_1 U14587 ( .A(n15289), .B(n15389), .C(n15373), .Y(n15149) );
  inv_1 U14588 ( .A(n15292), .Y(n15373) );
  nand2_1 U14589 ( .A(n15393), .B(n15444), .Y(n15292) );
  inv_1 U14590 ( .A(n15305), .Y(n15393) );
  nand2_1 U14591 ( .A(n23872), .B(n23895), .Y(n15305) );
  and3_1 U14592 ( .A(n15327), .B(n15454), .C(n15319), .X(n15289) );
  o21ai_0 U14593 ( .A1(n15019), .A2(n15107), .B1(n14965), .Y(n15451) );
  inv_1 U14594 ( .A(n14997), .Y(n14965) );
  nand2_1 U14595 ( .A(n15455), .B(n14964), .Y(n14997) );
  inv_1 U14596 ( .A(n15453), .Y(n15455) );
  nand2_1 U14597 ( .A(n15449), .B(n15448), .Y(n15453) );
  inv_1 U14598 ( .A(n15075), .Y(n15107) );
  nand3_1 U14599 ( .A(n15205), .B(n14851), .C(n15456), .Y(n15075) );
  nor3_1 U14600 ( .A(n15438), .B(n23871), .C(n23836), .Y(n15456) );
  inv_1 U14601 ( .A(n15259), .Y(n14851) );
  nand2_1 U14602 ( .A(n15359), .B(n15214), .Y(n15259) );
  nor2_1 U14603 ( .A(n15433), .B(n15304), .Y(n15214) );
  nor2_1 U14604 ( .A(n15457), .B(n23872), .Y(n15359) );
  and2_0 U14605 ( .A(n15319), .B(n15362), .X(n15205) );
  nor2_1 U14606 ( .A(n15187), .B(n24037), .Y(n15319) );
  nand2_1 U14607 ( .A(n23837), .B(n23893), .Y(n15187) );
  inv_1 U14608 ( .A(n15057), .Y(n15019) );
  nand3_1 U14609 ( .A(n14919), .B(n14920), .C(n15313), .Y(n15057) );
  inv_1 U14610 ( .A(n15258), .Y(n15313) );
  nand2_1 U14611 ( .A(n15454), .B(n23892), .Y(n15258) );
  nor2_1 U14612 ( .A(n15372), .B(n23895), .Y(n14919) );
  inv_1 U14613 ( .A(n23872), .Y(n15372) );
  or2_0 U14614 ( .A(n14943), .B(n14942), .X(n15450) );
  inv_1 U14615 ( .A(n14864), .Y(n14942) );
  nor2_1 U14616 ( .A(n15447), .B(n14859), .Y(n14864) );
  inv_1 U14617 ( .A(n14964), .Y(n14859) );
  nand3_1 U14618 ( .A(n15458), .B(n24051), .C(n15459), .Y(n14964) );
  nor2_1 U14619 ( .A(n15449), .B(inData[1]), .Y(n15447) );
  nand4_1 U14620 ( .A(n15327), .B(n15454), .C(n15389), .D(n15460), .Y(n14943)
         );
  nor2_1 U14621 ( .A(n14962), .B(n15365), .Y(n15460) );
  nand2_1 U14622 ( .A(n15243), .B(n23893), .Y(n15365) );
  inv_1 U14623 ( .A(n14982), .Y(n15243) );
  nand2_1 U14624 ( .A(n14873), .B(n10614), .Y(n14982) );
  nand2_1 U14625 ( .A(n14909), .B(n15444), .Y(n14962) );
  nor2_1 U14626 ( .A(n15398), .B(n15445), .Y(n15389) );
  inv_1 U14627 ( .A(n15430), .Y(n15327) );
  nand2_1 U14628 ( .A(n23873), .B(n23892), .Y(n15430) );
  o221ai_1 U14629 ( .A1(n15461), .A2(n11009), .B1(n15462), .B2(n10977), .C1(
        n15463), .Y(n10362) );
  nor2_1 U14630 ( .A(n14714), .B(n15464), .Y(n15463) );
  a21oi_1 U14631 ( .A1(n15465), .A2(n15466), .B1(n14710), .Y(n15464) );
  and4_1 U14632 ( .A(n15467), .B(n15468), .C(n11024), .D(n14735), .X(n15466)
         );
  nor3_1 U14633 ( .A(n15469), .B(n14831), .C(n14720), .Y(n15467) );
  nor4_1 U14634 ( .A(n15470), .B(n15471), .C(n15472), .D(n14820), .Y(n15465)
         );
  nand4_1 U14635 ( .A(n14716), .B(n10995), .C(n15473), .D(n15474), .Y(n14820)
         );
  and4_1 U14636 ( .A(n14790), .B(n14724), .C(n15475), .D(n15476), .X(n15474)
         );
  nand3_1 U14637 ( .A(n15477), .B(n15478), .C(n15479), .Y(n15470) );
  inv_1 U14638 ( .A(n10978), .Y(n14714) );
  nor4_1 U14639 ( .A(n15480), .B(n15481), .C(n15482), .D(n15483), .Y(n15462)
         );
  nor2_1 U14640 ( .A(n15484), .B(n15485), .Y(n15482) );
  nand4_1 U14641 ( .A(n15486), .B(n15487), .C(n15488), .D(n14833), .Y(n15480)
         );
  nor4_1 U14642 ( .A(n15489), .B(n15490), .C(n15491), .D(n15492), .Y(n15461)
         );
  inv_1 U14643 ( .A(n14738), .Y(n15491) );
  nand3_1 U14644 ( .A(n15493), .B(n15494), .C(n15495), .Y(n15490) );
  nand4_1 U14645 ( .A(n15496), .B(n14818), .C(n15497), .D(n15498), .Y(n15489)
         );
  inv_1 U14646 ( .A(n15499), .Y(n15496) );
  o211ai_1 U14647 ( .A1(n11009), .A2(n15500), .B1(n10978), .C1(n15501), .Y(
        n10361) );
  mux2i_1 U14648 ( .A0(n14784), .A1(n15502), .S(n15503), .Y(n15501) );
  nor4_1 U14649 ( .A(n15504), .B(n15505), .C(n15481), .D(n15506), .Y(n15503)
         );
  nand4_1 U14650 ( .A(n15507), .B(n14794), .C(n15508), .D(n11003), .Y(n15481)
         );
  nand3_1 U14651 ( .A(n15509), .B(n15510), .C(n15511), .Y(n15505) );
  nand4_1 U14652 ( .A(n11007), .B(n15512), .C(n15494), .D(n15513), .Y(n15504)
         );
  nor2_1 U14653 ( .A(n14811), .B(n14776), .Y(n15513) );
  nor3_1 U14654 ( .A(n14710), .B(n15514), .C(n10998), .Y(n15502) );
  nor4_1 U14655 ( .A(n15515), .B(n15516), .C(n15517), .D(n14783), .Y(n15500)
         );
  nand2_1 U14656 ( .A(n15518), .B(n15519), .Y(n14783) );
  inv_1 U14657 ( .A(n15472), .Y(n15518) );
  o221ai_1 U14658 ( .A1(n15520), .A2(n11009), .B1(n15521), .B2(n14710), .C1(
        n15522), .Y(n10360) );
  a21oi_1 U14659 ( .A1(n14784), .A2(n15523), .B1(n15524), .Y(n15522) );
  nand4_1 U14660 ( .A(n15525), .B(n15526), .C(n14826), .D(n15527), .Y(n15523)
         );
  nor3_1 U14661 ( .A(n15469), .B(n15528), .C(n15529), .Y(n15527) );
  inv_1 U14662 ( .A(n14733), .Y(n15525) );
  nand4_1 U14663 ( .A(n10995), .B(n15519), .C(n15530), .D(n15531), .Y(n14733)
         );
  and3_1 U14664 ( .A(n10994), .B(n15532), .C(n15508), .X(n15531) );
  nor4_1 U14665 ( .A(n15533), .B(n15534), .C(n15535), .D(n15536), .Y(n15521)
         );
  nand3_1 U14666 ( .A(n14778), .B(n15537), .C(n14791), .Y(n15534) );
  nand4_1 U14667 ( .A(n15538), .B(n15539), .C(n15540), .D(n14816), .Y(n15533)
         );
  inv_1 U14668 ( .A(n15541), .Y(n15539) );
  nor3_1 U14669 ( .A(n15542), .B(n14795), .C(n15543), .Y(n15520) );
  nand4_1 U14670 ( .A(n15544), .B(n14726), .C(n15545), .D(n15546), .Y(n14795)
         );
  inv_1 U14671 ( .A(n14825), .Y(n15544) );
  nand3_1 U14672 ( .A(n15497), .B(n11003), .C(n14734), .Y(n15542) );
  nand4_1 U14673 ( .A(n15547), .B(n15548), .C(n14769), .D(n10978), .Y(n10359)
         );
  nand2_1 U14674 ( .A(n15524), .B(n15452), .Y(n10978) );
  inv_1 U14675 ( .A(n15360), .Y(n15452) );
  o21ai_0 U14676 ( .A1(n15549), .A2(n15550), .B1(n14302), .Y(n15548) );
  nand4_1 U14677 ( .A(n15526), .B(n15551), .C(n15552), .D(n15553), .Y(n15550)
         );
  nor2_1 U14678 ( .A(n15554), .B(n15555), .Y(n15553) );
  nand4_1 U14679 ( .A(n15509), .B(n10995), .C(n15556), .D(n15557), .Y(n15549)
         );
  nor2_1 U14680 ( .A(n11011), .B(n15558), .Y(n15556) );
  mux2i_1 U14681 ( .A0(n10980), .A1(n15559), .S(n15560), .Y(n15547) );
  nor4_1 U14682 ( .A(n15561), .B(n15562), .C(n15563), .D(n15564), .Y(n15560)
         );
  nand2_1 U14683 ( .A(n14818), .B(n14808), .Y(n15562) );
  nand4_1 U14684 ( .A(n15476), .B(n15565), .C(n14765), .D(n10991), .Y(n15561)
         );
  nor4_1 U14685 ( .A(n15566), .B(n15567), .C(n10998), .D(n15568), .Y(n15559)
         );
  or3_1 U14686 ( .A(n10977), .B(n15569), .C(n15570), .X(n15567) );
  nand3_1 U14687 ( .A(n15519), .B(n15571), .C(n15572), .Y(n15566) );
  and3_1 U14688 ( .A(n14723), .B(n15573), .C(n14821), .X(n15572) );
  o21ai_0 U14689 ( .A1(n15574), .A2(n11009), .B1(n15575), .Y(n10358) );
  mux2i_1 U14690 ( .A0(n14784), .A1(n15576), .S(n15577), .Y(n15575) );
  nor4_1 U14691 ( .A(n15578), .B(n15579), .C(n15580), .D(n15581), .Y(n15577)
         );
  nand2_1 U14692 ( .A(n15582), .B(n15583), .Y(n15579) );
  inv_1 U14693 ( .A(n15471), .Y(n15583) );
  nand4_1 U14694 ( .A(n14734), .B(n14836), .C(n15571), .D(n15584), .Y(n15471)
         );
  nand4_1 U14695 ( .A(n15497), .B(n15565), .C(n14821), .D(n15495), .Y(n15578)
         );
  nor4_1 U14696 ( .A(n15585), .B(n15586), .C(n15587), .D(n15588), .Y(n15576)
         );
  or3_1 U14697 ( .A(n15589), .B(n15590), .C(n15591), .X(n15586) );
  nand4_1 U14698 ( .A(n15592), .B(n14764), .C(n14779), .D(n15593), .Y(n15585)
         );
  nor3_1 U14699 ( .A(n15594), .B(n11020), .C(n14720), .Y(n15593) );
  inv_1 U14700 ( .A(n15595), .Y(n14720) );
  nor4_1 U14701 ( .A(n15596), .B(n15499), .C(n14729), .D(n14732), .Y(n15574)
         );
  nand4_1 U14702 ( .A(n15545), .B(n11007), .C(n15498), .D(n15597), .Y(n14732)
         );
  nor3_1 U14703 ( .A(n15569), .B(n15598), .C(n15599), .Y(n15597) );
  nand3_1 U14704 ( .A(n14791), .B(n10990), .C(n11004), .Y(n14729) );
  inv_1 U14705 ( .A(n15600), .Y(n11004) );
  nand3_1 U14706 ( .A(n15519), .B(n15573), .C(n10989), .Y(n15499) );
  nand4_1 U14707 ( .A(n15509), .B(n14807), .C(n14778), .D(n14754), .Y(n15596)
         );
  o21ai_0 U14708 ( .A1(n15601), .A2(n14710), .B1(n15602), .Y(n10357) );
  mux2i_1 U14709 ( .A0(n14784), .A1(n15603), .S(n15604), .Y(n15602) );
  nor4_1 U14710 ( .A(n15605), .B(n14823), .C(n15606), .D(n14777), .Y(n15604)
         );
  inv_1 U14711 ( .A(n11007), .Y(n15606) );
  nand2_1 U14712 ( .A(n15607), .B(n15538), .Y(n15605) );
  and3_1 U14713 ( .A(n15584), .B(n15608), .C(n15609), .X(n15538) );
  nor4_1 U14714 ( .A(n15610), .B(n15611), .C(n15612), .D(n14782), .Y(n15603)
         );
  nand3_1 U14715 ( .A(n14302), .B(n15613), .C(n14724), .Y(n15611) );
  nand3_1 U14716 ( .A(n15601), .B(n15582), .C(n15614), .Y(n15610) );
  nor3_1 U14717 ( .A(n15541), .B(n15615), .C(n15543), .Y(n15614) );
  nand4_1 U14718 ( .A(n15486), .B(n15557), .C(n14836), .D(n15616), .Y(n15543)
         );
  nor4_1 U14719 ( .A(n15617), .B(n14832), .C(n15618), .D(n15619), .Y(n15616)
         );
  inv_1 U14720 ( .A(n10990), .Y(n14832) );
  nand4_1 U14721 ( .A(n14808), .B(n15476), .C(n15620), .D(n15621), .Y(n15541)
         );
  and3_1 U14722 ( .A(n14835), .B(n15488), .C(n14740), .X(n15621) );
  and3_1 U14723 ( .A(n15622), .B(n15508), .C(n14838), .X(n15582) );
  and4_1 U14724 ( .A(n15623), .B(n15540), .C(n15624), .D(n15625), .X(n15601)
         );
  and4_1 U14725 ( .A(n15626), .B(n15498), .C(n14791), .D(n15475), .X(n15625)
         );
  and4_1 U14726 ( .A(n14790), .B(n15493), .C(n11003), .D(n14737), .X(n15626)
         );
  nor3_1 U14727 ( .A(n14804), .B(n15627), .C(n15628), .Y(n15624) );
  nand3_1 U14728 ( .A(n15519), .B(n15629), .C(n15477), .Y(n14804) );
  inv_1 U14729 ( .A(n15630), .Y(n15477) );
  nor2_1 U14730 ( .A(n14776), .B(n15589), .Y(n15623) );
  inv_1 U14731 ( .A(n15497), .Y(n14776) );
  o22ai_1 U14732 ( .A1(n10924), .A2(n11014), .B1(n11703), .B2(n15631), .Y(
        n10356) );
  xor2_1 U14733 ( .A(outData[27]), .B(n11497), .X(n15631) );
  inv_1 U14734 ( .A(n12587), .Y(n11014) );
  nand4_1 U14735 ( .A(n15632), .B(n15633), .C(n15634), .D(n14768), .Y(n10355)
         );
  o21ai_0 U14736 ( .A1(n15635), .A2(n15636), .B1(n14784), .Y(n15634) );
  or4_1 U14737 ( .A(n15555), .B(n15472), .C(n15637), .D(n15638), .X(n15636) );
  nand3_1 U14738 ( .A(n15530), .B(n11024), .C(n15498), .Y(n15638) );
  inv_1 U14739 ( .A(n15568), .Y(n15530) );
  nand3_1 U14740 ( .A(n14806), .B(n14790), .C(n14838), .Y(n15568) );
  nand4_1 U14741 ( .A(n11026), .B(n15639), .C(n15557), .D(n14725), .Y(n15472)
         );
  nand3_1 U14742 ( .A(n14736), .B(n15493), .C(n14763), .Y(n15555) );
  nand4_1 U14743 ( .A(n14809), .B(n11007), .C(n15592), .D(n15640), .Y(n15635)
         );
  nor3_1 U14744 ( .A(n15558), .B(n14721), .C(n14722), .Y(n15640) );
  inv_1 U14745 ( .A(n15641), .Y(n14722) );
  inv_1 U14746 ( .A(n15642), .Y(n15558) );
  nand2_1 U14747 ( .A(n10980), .B(n15643), .Y(n15633) );
  nand4_1 U14748 ( .A(n14734), .B(n10994), .C(n15644), .D(n15645), .Y(n15643)
         );
  nor4_1 U14749 ( .A(n14744), .B(n14796), .C(n14805), .D(n15591), .Y(n15645)
         );
  nand3_1 U14750 ( .A(n15646), .B(n15647), .C(n14726), .Y(n15591) );
  nand3_1 U14751 ( .A(n15620), .B(n15648), .C(n15649), .Y(n14805) );
  inv_1 U14752 ( .A(n15628), .Y(n15649) );
  nand4_1 U14753 ( .A(n14758), .B(n15650), .C(n15651), .D(n14765), .Y(n15628)
         );
  nor3_1 U14754 ( .A(n15652), .B(n15653), .C(n15590), .Y(n15620) );
  nand3_1 U14755 ( .A(n15487), .B(n15512), .C(n15571), .Y(n14744) );
  nor3_1 U14756 ( .A(n14757), .B(n14750), .C(n15529), .Y(n15644) );
  inv_1 U14757 ( .A(n14778), .Y(n14750) );
  o21ai_0 U14758 ( .A1(n15654), .A2(n15655), .B1(n14302), .Y(n15632) );
  nand4_1 U14759 ( .A(n14771), .B(n15551), .C(n14818), .D(n15656), .Y(n15655)
         );
  and3_1 U14760 ( .A(n15486), .B(n15595), .C(n14727), .X(n15656) );
  and4_1 U14761 ( .A(n10990), .B(n14724), .C(n15479), .D(n15657), .X(n14771)
         );
  and4_1 U14762 ( .A(n10991), .B(n11003), .C(n14764), .D(n15495), .X(n15657)
         );
  and4_1 U14763 ( .A(n15658), .B(n15510), .C(n10992), .D(n15659), .X(n15479)
         );
  nand4_1 U14764 ( .A(n14835), .B(n14837), .C(n15608), .D(n15660), .Y(n15654)
         );
  and4_1 U14765 ( .A(n14833), .B(n15488), .C(n14754), .D(n14821), .X(n15660)
         );
  o221ai_1 U14766 ( .A1(n11009), .A2(n15661), .B1(n15662), .B2(n14710), .C1(
        n15663), .Y(n10354) );
  o22ai_1 U14767 ( .A1(n14784), .A2(n15664), .B1(n15665), .B2(n15666), .Y(
        n15663) );
  nand4_1 U14768 ( .A(n15607), .B(n14760), .C(n15667), .D(n15668), .Y(n15666)
         );
  nor3_1 U14769 ( .A(n11029), .B(n15669), .C(n15670), .Y(n15668) );
  nand3_1 U14770 ( .A(n15508), .B(n15592), .C(n15509), .Y(n11029) );
  and3_1 U14771 ( .A(n11001), .B(n14835), .C(n15671), .X(n14760) );
  and3_1 U14772 ( .A(n14779), .B(n15648), .C(n14821), .X(n15671) );
  and3_1 U14773 ( .A(n14778), .B(n15532), .C(n10995), .X(n15607) );
  nand4_1 U14774 ( .A(n14791), .B(n10992), .C(n15622), .D(n15672), .Y(n15665)
         );
  and4_1 U14775 ( .A(n15651), .B(n15488), .C(n14754), .D(n14738), .X(n15672)
         );
  nor4_1 U14776 ( .A(n15673), .B(n15674), .C(n14796), .D(n15588), .Y(n15662)
         );
  nand3_1 U14777 ( .A(n14806), .B(n15659), .C(n15675), .Y(n15588) );
  or3_1 U14778 ( .A(n10986), .B(n15516), .C(n15627), .X(n15674) );
  nand4_1 U14779 ( .A(n11016), .B(n15584), .C(n15676), .D(n14725), .Y(n15673)
         );
  nor2_1 U14780 ( .A(n15617), .B(n15677), .Y(n15676) );
  inv_1 U14781 ( .A(n10991), .Y(n15617) );
  inv_1 U14782 ( .A(n14824), .Y(n11016) );
  nand3_1 U14783 ( .A(n15678), .B(n15507), .C(n15679), .Y(n14824) );
  and3_1 U14784 ( .A(n14728), .B(n15546), .C(n15545), .X(n15679) );
  inv_1 U14785 ( .A(n15680), .Y(n15507) );
  nor4_1 U14786 ( .A(n14812), .B(n14759), .C(n14825), .D(n15563), .Y(n15661)
         );
  nand2_1 U14787 ( .A(n14809), .B(n10994), .Y(n15563) );
  o211ai_1 U14788 ( .A1(n15681), .A2(n10977), .B1(n15682), .C1(n15683), .Y(
        n10353) );
  o21ai_0 U14789 ( .A1(n15684), .A2(n15685), .B1(n14302), .Y(n15683) );
  nand4_1 U14790 ( .A(n15686), .B(n15609), .C(n11000), .D(n15551), .Y(n15685)
         );
  nor3_1 U14791 ( .A(n15492), .B(n14811), .C(n14777), .Y(n11000) );
  inv_1 U14792 ( .A(n14740), .Y(n15492) );
  and4_1 U14793 ( .A(n14794), .B(n11026), .C(n14821), .D(n15494), .X(n15609)
         );
  nand4_1 U14794 ( .A(n15510), .B(n14725), .C(n15648), .D(n14790), .Y(n15684)
         );
  o22ai_1 U14795 ( .A1(n10980), .A2(n15664), .B1(n15687), .B2(n15688), .Y(
        n15682) );
  nand4_1 U14796 ( .A(n15689), .B(n15511), .C(n15667), .D(n15690), .Y(n15688)
         );
  nor3_1 U14797 ( .A(n15590), .B(n15680), .C(n10985), .Y(n15690) );
  nor3_1 U14798 ( .A(n14831), .B(n11011), .C(n15664), .Y(n15667) );
  inv_1 U14799 ( .A(n14737), .Y(n11011) );
  inv_1 U14800 ( .A(n15564), .Y(n15689) );
  nand4_1 U14801 ( .A(n10990), .B(n11007), .C(n15691), .D(n15692), .Y(n15564)
         );
  nor4_1 U14802 ( .A(n15693), .B(n15599), .C(n15630), .D(n14797), .Y(n15692)
         );
  nand3_1 U14803 ( .A(n15498), .B(n15629), .C(n15473), .Y(n14797) );
  inv_1 U14804 ( .A(n15627), .Y(n15473) );
  inv_1 U14805 ( .A(n15486), .Y(n15599) );
  nor3_1 U14806 ( .A(n11010), .B(n15653), .C(n15652), .Y(n15691) );
  inv_1 U14807 ( .A(n14753), .Y(n15652) );
  inv_1 U14808 ( .A(n15694), .Y(n15653) );
  inv_1 U14809 ( .A(n15512), .Y(n11010) );
  nand4_1 U14810 ( .A(n14764), .B(n15493), .C(n14837), .D(n15695), .Y(n15687)
         );
  nor3_1 U14811 ( .A(n15696), .B(n14757), .C(n15697), .Y(n15695) );
  inv_1 U14812 ( .A(n15476), .Y(n15696) );
  inv_1 U14813 ( .A(n14768), .Y(n15664) );
  nand2_1 U14814 ( .A(n15524), .B(n15360), .Y(n14768) );
  nand3_1 U14815 ( .A(n14920), .B(n15410), .C(n14909), .Y(n15360) );
  nor2_1 U14816 ( .A(n23872), .B(n23895), .Y(n14909) );
  inv_1 U14817 ( .A(n15438), .Y(n15410) );
  nand2_1 U14818 ( .A(n15454), .B(n15184), .Y(n15438) );
  inv_1 U14819 ( .A(n14890), .Y(n15454) );
  nand2_1 U14820 ( .A(n15435), .B(n10774), .Y(n14890) );
  and3_1 U14821 ( .A(n15357), .B(n15444), .C(n12462), .X(n14920) );
  nor2_1 U14822 ( .A(n14873), .B(n23837), .Y(n12462) );
  nor2_1 U14823 ( .A(n15433), .B(n23894), .Y(n15444) );
  inv_1 U14824 ( .A(n24036), .Y(n15433) );
  nor3_1 U14825 ( .A(n23836), .B(n23871), .C(n15370), .Y(n15357) );
  nand2_1 U14826 ( .A(n15311), .B(n15362), .Y(n15370) );
  inv_1 U14827 ( .A(n14710), .Y(n10980) );
  nor4_1 U14828 ( .A(n15698), .B(n15699), .C(n15670), .D(n15637), .Y(n15681)
         );
  nand4_1 U14829 ( .A(n14728), .B(n11030), .C(n14826), .D(n15700), .Y(n15637)
         );
  and4_1 U14830 ( .A(n15573), .B(n14723), .C(n14836), .D(n10995), .X(n15700)
         );
  and2_0 U14831 ( .A(n15509), .B(n15622), .X(n14826) );
  inv_1 U14832 ( .A(n15658), .Y(n15670) );
  nand3_1 U14833 ( .A(n15519), .B(n14806), .C(n15557), .Y(n15699) );
  nand4_1 U14834 ( .A(n14754), .B(n11003), .C(n14809), .D(n15701), .Y(n15698)
         );
  and2_0 U14835 ( .A(n15545), .B(n15508), .X(n15701) );
  o211ai_1 U14836 ( .A1(n15702), .A2(n11009), .B1(n14769), .C1(n15703), .Y(
        n10352) );
  mux2i_1 U14837 ( .A0(n14784), .A1(n15704), .S(n15705), .Y(n15703) );
  nor4_1 U14838 ( .A(n15706), .B(n15707), .C(n15598), .D(n14777), .Y(n15705)
         );
  inv_1 U14839 ( .A(n14734), .Y(n14777) );
  inv_1 U14840 ( .A(n15557), .Y(n15598) );
  nand3_1 U14841 ( .A(n11005), .B(n14833), .C(n14725), .Y(n15707) );
  nand4_1 U14842 ( .A(n15708), .B(n15468), .C(n10989), .D(n10995), .Y(n15706)
         );
  inv_1 U14843 ( .A(n15506), .Y(n15708) );
  nand4_1 U14844 ( .A(n15622), .B(n14791), .C(n14836), .D(n15709), .Y(n15506)
         );
  and3_1 U14845 ( .A(n14838), .B(n14746), .C(n11015), .X(n15709) );
  inv_1 U14846 ( .A(n15710), .Y(n14838) );
  o21ai_0 U14847 ( .A1(n10987), .A2(n10988), .B1(n15711), .Y(n15710) );
  nand4_1 U14848 ( .A(n15712), .B(n15713), .C(n15714), .D(n15715), .Y(n15711)
         );
  nand4_1 U14849 ( .A(n15716), .B(n15715), .C(n15717), .D(n15718), .Y(n10988)
         );
  inv_1 U14850 ( .A(n15719), .Y(n10987) );
  nor4_1 U14851 ( .A(n15720), .B(n15721), .C(n15587), .D(n15722), .Y(n15704)
         );
  nand2_1 U14852 ( .A(n14818), .B(n15723), .Y(n15722) );
  inv_1 U14853 ( .A(n14796), .Y(n15723) );
  nand2_1 U14854 ( .A(n15475), .B(n15494), .Y(n14796) );
  and2_0 U14855 ( .A(n14741), .B(n15532), .X(n14818) );
  nand4_1 U14856 ( .A(n15526), .B(n15642), .C(n15724), .D(n15725), .Y(n15587)
         );
  and4_1 U14857 ( .A(n14737), .B(n15726), .C(n14724), .D(n11025), .X(n15725)
         );
  nor2_1 U14858 ( .A(n10998), .B(n14710), .Y(n15724) );
  nand2_1 U14859 ( .A(n15727), .B(n15613), .Y(n10998) );
  nand4_1 U14860 ( .A(n15728), .B(n15729), .C(n15730), .D(n15731), .Y(n15613)
         );
  and4_1 U14861 ( .A(n15732), .B(n15727), .C(n14765), .D(n14753), .X(n15731)
         );
  nand4_1 U14862 ( .A(n15713), .B(n15733), .C(n15734), .D(n15735), .Y(n14753)
         );
  o21ai_0 U14863 ( .A1(n15736), .A2(n15737), .B1(n15735), .Y(n14765) );
  and3_1 U14864 ( .A(n15738), .B(n15717), .C(n15739), .X(n15737) );
  nor4_1 U14865 ( .A(n24051), .B(n15740), .C(n15741), .D(n11133), .Y(n15736)
         );
  nor2_1 U14866 ( .A(n11020), .B(n14811), .Y(n15732) );
  inv_1 U14867 ( .A(n15537), .Y(n14811) );
  inv_1 U14868 ( .A(n15629), .Y(n11020) );
  nand4_1 U14869 ( .A(n15742), .B(n15743), .C(n15744), .D(n15745), .Y(n15629)
         );
  nor4_1 U14870 ( .A(n15669), .B(n14759), .C(n10986), .D(n14789), .Y(n15730)
         );
  nand4_1 U14871 ( .A(n15552), .B(n11015), .C(n15540), .D(n15746), .Y(n14789)
         );
  and4_1 U14872 ( .A(n11007), .B(n14807), .C(n10994), .D(n15622), .X(n15746)
         );
  nand4_1 U14873 ( .A(n15747), .B(n15738), .C(n15748), .D(n15717), .Y(n15622)
         );
  and3_1 U14874 ( .A(n14716), .B(n14762), .C(n15511), .X(n15540) );
  inv_1 U14875 ( .A(n15749), .Y(n15511) );
  nor4_1 U14876 ( .A(n14721), .B(n15697), .C(n15619), .D(n15612), .Y(n11015)
         );
  inv_1 U14877 ( .A(n14763), .Y(n15619) );
  inv_1 U14878 ( .A(n15608), .Y(n15697) );
  nand2_1 U14879 ( .A(n15750), .B(n15751), .Y(n15608) );
  inv_1 U14880 ( .A(n15584), .Y(n14721) );
  nand4_1 U14881 ( .A(n15752), .B(n15753), .C(n15754), .D(n15755), .Y(n15584)
         );
  inv_1 U14882 ( .A(n15516), .Y(n15552) );
  nand2_1 U14883 ( .A(n14816), .B(n14833), .Y(n15516) );
  inv_1 U14884 ( .A(n15589), .Y(n14816) );
  nand4_1 U14885 ( .A(n15486), .B(n15476), .C(n15639), .D(n15756), .Y(n10986)
         );
  and4_1 U14886 ( .A(n15694), .B(n15498), .C(n15519), .D(n15557), .X(n15756)
         );
  nand4_1 U14887 ( .A(n15757), .B(n15758), .C(n15742), .D(n15745), .Y(n15557)
         );
  nand4_1 U14888 ( .A(n15757), .B(n15733), .C(n15734), .D(n15744), .Y(n15694)
         );
  nand4_1 U14889 ( .A(n15759), .B(n15760), .C(n15761), .D(n15762), .Y(n15486)
         );
  nand3_1 U14890 ( .A(n15497), .B(n14836), .C(n15510), .Y(n14759) );
  nand4_1 U14891 ( .A(n15763), .B(n15754), .C(n15755), .D(n15764), .Y(n14836)
         );
  nand3_1 U14892 ( .A(n15765), .B(n15761), .C(n15766), .Y(n15497) );
  nor4_1 U14893 ( .A(n15767), .B(n15627), .C(n15570), .D(n15517), .Y(n15729)
         );
  nand2_1 U14894 ( .A(n15768), .B(n15769), .Y(n15517) );
  nor4_1 U14895 ( .A(n15770), .B(n15771), .C(n14831), .D(n14812), .Y(n15769)
         );
  inv_1 U14896 ( .A(n15573), .Y(n14812) );
  nand3_1 U14897 ( .A(n15772), .B(n15752), .C(n15757), .Y(n15573) );
  inv_1 U14898 ( .A(n14754), .Y(n15771) );
  nand3_1 U14899 ( .A(n15739), .B(n15745), .C(n15773), .Y(n14754) );
  nand4_1 U14900 ( .A(n14790), .B(n14736), .C(n14764), .D(n15532), .Y(n15770)
         );
  nor4_1 U14901 ( .A(n15774), .B(n15615), .C(n15483), .D(n14823), .Y(n15768)
         );
  nand4_1 U14902 ( .A(n14778), .B(n15592), .C(n14821), .D(n15775), .Y(n15483)
         );
  and4_1 U14903 ( .A(n10991), .B(n15648), .C(n14809), .D(n15546), .X(n15775)
         );
  nand4_1 U14904 ( .A(n15738), .B(n15757), .C(n15713), .D(n15717), .Y(n14821)
         );
  nand3_1 U14905 ( .A(n15776), .B(n15777), .C(n15772), .Y(n14778) );
  nand4_1 U14906 ( .A(n15468), .B(n10990), .C(n14724), .D(n15659), .Y(n15774)
         );
  nand4_1 U14907 ( .A(n15778), .B(n15752), .C(n15762), .D(n15779), .Y(n14724)
         );
  nor3_1 U14908 ( .A(n14751), .B(n11021), .C(n15677), .Y(n15468) );
  inv_1 U14909 ( .A(n14837), .Y(n15677) );
  nand4_1 U14910 ( .A(n15748), .B(n15735), .C(n15776), .D(n15745), .Y(n14837)
         );
  inv_1 U14911 ( .A(n14723), .Y(n11021) );
  inv_1 U14912 ( .A(n15780), .Y(n14751) );
  nand4_1 U14913 ( .A(n15478), .B(n15781), .C(n15782), .D(n15783), .Y(n15570)
         );
  nor4_1 U14914 ( .A(n15784), .B(n15785), .C(n15528), .D(n15618), .Y(n15783)
         );
  inv_1 U14915 ( .A(n14725), .Y(n15618) );
  nand3_1 U14916 ( .A(n15772), .B(n15786), .C(n15747), .Y(n14725) );
  inv_1 U14917 ( .A(n10992), .Y(n15528) );
  nand2_1 U14918 ( .A(n15545), .B(n11003), .Y(n15785) );
  and3_1 U14919 ( .A(n14758), .B(n15508), .C(n14740), .X(n15782) );
  nand2_1 U14920 ( .A(n15458), .B(n15761), .Y(n14740) );
  nand2_1 U14921 ( .A(n15787), .B(n15748), .Y(n14758) );
  inv_1 U14922 ( .A(n10985), .Y(n15781) );
  nand4_1 U14923 ( .A(n14835), .B(n15475), .C(n14791), .D(n14779), .Y(n10985)
         );
  nand4_1 U14924 ( .A(n15788), .B(n15712), .C(n15789), .D(n15748), .Y(n15475)
         );
  nand2_1 U14925 ( .A(n15790), .B(n15791), .Y(n15627) );
  nand4_1 U14926 ( .A(n15757), .B(n15734), .C(n15758), .D(n15792), .Y(n15791)
         );
  nand3_1 U14927 ( .A(n15772), .B(n15777), .C(n15712), .Y(n15790) );
  inv_1 U14928 ( .A(n14808), .Y(n15767) );
  nor4_1 U14929 ( .A(n14757), .B(n15793), .C(n15794), .D(n11012), .Y(n14808)
         );
  inv_1 U14930 ( .A(n15726), .Y(n11012) );
  and3_1 U14931 ( .A(n15713), .B(n15714), .C(n15773), .X(n14757) );
  nor3_1 U14932 ( .A(n24051), .B(n24052), .C(n15795), .Y(n15713) );
  nor4_1 U14933 ( .A(n15630), .B(n15600), .C(n15554), .D(n15796), .Y(n15728)
         );
  nand2_1 U14934 ( .A(n14746), .B(n14726), .Y(n15554) );
  inv_1 U14935 ( .A(n15536), .Y(n14746) );
  nand2_1 U14936 ( .A(n15658), .B(n14834), .Y(n15536) );
  nand4_1 U14937 ( .A(n15797), .B(n15798), .C(n15799), .D(n15800), .Y(n15658)
         );
  nor2_1 U14938 ( .A(n11400), .B(n15801), .Y(n15800) );
  nand4_1 U14939 ( .A(n15488), .B(n15493), .C(n15651), .D(n15494), .Y(n15600)
         );
  nand2_1 U14940 ( .A(n15802), .B(n15764), .Y(n15493) );
  nand3_1 U14941 ( .A(n15789), .B(n15764), .C(n15803), .Y(n15488) );
  inv_1 U14942 ( .A(n14823), .Y(n15526) );
  nand2_1 U14943 ( .A(n14738), .B(n15487), .Y(n14823) );
  nand3_1 U14944 ( .A(n14735), .B(n14727), .C(n14761), .Y(n15721) );
  and3_1 U14945 ( .A(n15476), .B(n11006), .C(n14817), .X(n14761) );
  nand2_1 U14946 ( .A(n15804), .B(n15792), .Y(n15476) );
  nand4_1 U14947 ( .A(n10994), .B(n15508), .C(n15565), .D(n15805), .Y(n15720)
         );
  and3_1 U14948 ( .A(n11023), .B(n14752), .C(n15537), .X(n15805) );
  nand3_1 U14949 ( .A(n15806), .B(n15742), .C(n15807), .Y(n15508) );
  inv_1 U14950 ( .A(n10977), .Y(n14784) );
  nor4_1 U14951 ( .A(n15808), .B(n15809), .C(n15693), .D(n15569), .Y(n15702)
         );
  inv_1 U14952 ( .A(n15639), .Y(n15569) );
  nand2_1 U14953 ( .A(n15810), .B(n15715), .Y(n15639) );
  inv_1 U14954 ( .A(n15592), .Y(n15693) );
  nand2_1 U14955 ( .A(n15804), .B(n15752), .Y(n15592) );
  and3_1 U14956 ( .A(n15758), .B(n15714), .C(n15757), .X(n15804) );
  nand3_1 U14957 ( .A(n15659), .B(n15651), .C(n10990), .Y(n15809) );
  nand3_1 U14958 ( .A(n15715), .B(n15799), .C(n15772), .Y(n10990) );
  nand2_1 U14959 ( .A(n15802), .B(n15761), .Y(n15651) );
  and3_1 U14960 ( .A(n15760), .B(n15762), .C(n15712), .X(n15802) );
  nand4_1 U14961 ( .A(n15715), .B(n15718), .C(n15734), .D(n15811), .Y(n15659)
         );
  nor2_1 U14962 ( .A(n11133), .B(n15812), .Y(n15811) );
  or4_1 U14963 ( .A(n15813), .B(n15581), .C(n15535), .D(n15669), .X(n15808) );
  inv_1 U14964 ( .A(n11026), .Y(n15669) );
  nand4_1 U14965 ( .A(n15719), .B(n15758), .C(n15715), .D(n15717), .Y(n11026)
         );
  inv_1 U14966 ( .A(n15510), .Y(n15535) );
  nand4_1 U14967 ( .A(n14781), .B(n15806), .C(n15761), .D(n15742), .Y(n15510)
         );
  nand3_1 U14968 ( .A(n14835), .B(n15512), .C(n14794), .Y(n15581) );
  nand4_1 U14969 ( .A(n15789), .B(n12916), .C(n15814), .D(n15815), .Y(n14835)
         );
  and2_0 U14970 ( .A(n15764), .B(n15816), .X(n15814) );
  o221ai_1 U14971 ( .A1(n15817), .A2(n10977), .B1(n15818), .B2(n11009), .C1(
        n15819), .Y(n10351) );
  nor3_1 U14972 ( .A(n15820), .B(n15524), .C(n15821), .Y(n15819) );
  inv_1 U14973 ( .A(n14769), .Y(n15821) );
  nand2_1 U14974 ( .A(n14831), .B(n14302), .Y(n14769) );
  and4_1 U14975 ( .A(n15758), .B(n15786), .C(n15735), .D(n15714), .X(n14831)
         );
  nor2_1 U14976 ( .A(n15727), .B(n11009), .Y(n15524) );
  nand2_1 U14977 ( .A(n15799), .B(n15822), .Y(n15727) );
  a21oi_1 U14978 ( .A1(n15823), .A2(n15824), .B1(n14710), .Y(n15820) );
  nand2_1 U14979 ( .A(n12699), .B(n14302), .Y(n14710) );
  nor4_1 U14980 ( .A(n15825), .B(n15612), .C(n15794), .D(n15793), .Y(n15824)
         );
  inv_1 U14981 ( .A(n11025), .Y(n15793) );
  nand4_1 U14982 ( .A(n15786), .B(n15739), .C(n15735), .D(n15745), .Y(n11025)
         );
  inv_1 U14983 ( .A(n15646), .Y(n15794) );
  nand4_1 U14984 ( .A(n15747), .B(n15738), .C(n15789), .D(n15739), .Y(n15646)
         );
  inv_1 U14985 ( .A(n14806), .Y(n15612) );
  nand4_1 U14986 ( .A(n15815), .B(n15761), .C(n15826), .D(n15816), .Y(n14806)
         );
  nor2_1 U14987 ( .A(n15827), .B(n11442), .Y(n15826) );
  nand4_1 U14988 ( .A(n15545), .B(n15546), .C(n15487), .D(n15726), .Y(n15825)
         );
  nand4_1 U14989 ( .A(n15757), .B(n15744), .C(n15776), .D(n15717), .Y(n15726)
         );
  nand2_1 U14990 ( .A(n15828), .B(n15829), .Y(n15487) );
  nand3_1 U14991 ( .A(n15830), .B(n15779), .C(n12916), .Y(n15546) );
  nand2_1 U14992 ( .A(n15831), .B(n15719), .Y(n15545) );
  nor4_1 U14993 ( .A(n15832), .B(n15813), .C(n15749), .D(n15630), .Y(n15823)
         );
  nand3_1 U14994 ( .A(n11006), .B(n15647), .C(n14752), .Y(n15630) );
  nand3_1 U14995 ( .A(n15739), .B(n15833), .C(n15719), .Y(n14752) );
  nand3_1 U14996 ( .A(n15772), .B(n15799), .C(n15747), .Y(n15647) );
  and2_0 U14997 ( .A(n15748), .B(n15714), .X(n15772) );
  nand2_1 U14998 ( .A(n15788), .B(n15810), .Y(n11006) );
  and3_1 U14999 ( .A(n15789), .B(n15744), .C(n15712), .X(n15810) );
  nand2_1 U15000 ( .A(n15678), .B(n14741), .Y(n15749) );
  nand3_1 U15001 ( .A(n15834), .B(n15743), .C(n15763), .Y(n14741) );
  and3_1 U15002 ( .A(n15595), .B(n15641), .C(n15571), .X(n15678) );
  nand2_1 U15003 ( .A(n14781), .B(n15830), .Y(n15571) );
  and3_1 U15004 ( .A(n15835), .B(n15836), .C(n15834), .X(n15830) );
  nand3_1 U15005 ( .A(n15834), .B(n15755), .C(n15733), .Y(n15641) );
  nand3_1 U15006 ( .A(n15816), .B(n15743), .C(n15778), .Y(n15595) );
  nand4_1 U15007 ( .A(n14764), .B(n11007), .C(n14790), .D(n15837), .Y(n15813)
         );
  nor3_1 U15008 ( .A(n15580), .B(n15529), .C(n15838), .Y(n15837) );
  inv_1 U15009 ( .A(n15509), .Y(n15838) );
  nand2_1 U15010 ( .A(n12916), .B(n15750), .Y(n15509) );
  and3_1 U15011 ( .A(n15753), .B(n15816), .C(n15760), .X(n15750) );
  inv_1 U15012 ( .A(n14779), .Y(n15529) );
  nand4_1 U15013 ( .A(n15792), .B(n15798), .C(n15761), .D(n15839), .Y(n14779)
         );
  nor2_1 U15014 ( .A(n11211), .B(n15801), .Y(n15839) );
  nand3_1 U15015 ( .A(n15648), .B(n14736), .C(n14809), .Y(n15580) );
  nand2_1 U15016 ( .A(n15787), .B(n15744), .Y(n14809) );
  and3_1 U15017 ( .A(n15786), .B(n15743), .C(n15734), .X(n15787) );
  nand4_1 U15018 ( .A(n15719), .B(n15744), .C(n15777), .D(n15717), .Y(n14736)
         );
  nand4_1 U15019 ( .A(n15734), .B(n15758), .C(n15792), .D(n15715), .Y(n15648)
         );
  nor3_1 U15020 ( .A(n24051), .B(n24055), .C(n10832), .Y(n15758) );
  nand2_1 U15021 ( .A(n15840), .B(n15799), .Y(n14790) );
  and2_0 U15022 ( .A(n15836), .B(n11314), .X(n15799) );
  nand4_1 U15023 ( .A(n15765), .B(n15806), .C(n15753), .D(n15755), .Y(n11007)
         );
  nand4_1 U15024 ( .A(n15738), .B(n15789), .C(n15748), .D(n15735), .Y(n14764)
         );
  nand3_1 U15025 ( .A(n15478), .B(n15498), .C(n14716), .Y(n15832) );
  inv_1 U15026 ( .A(n15515), .Y(n14716) );
  nand2_1 U15027 ( .A(n15642), .B(n15565), .Y(n15515) );
  nand4_1 U15028 ( .A(n15788), .B(n15733), .C(n15806), .D(n15829), .Y(n15565)
         );
  nand2_1 U15029 ( .A(n15828), .B(n15841), .Y(n15642) );
  and3_1 U15030 ( .A(n15734), .B(n15755), .C(n15738), .X(n15828) );
  nand4_1 U15031 ( .A(n15738), .B(n14781), .C(n15806), .D(n15764), .Y(n15498)
         );
  inv_1 U15032 ( .A(n15590), .Y(n15478) );
  nand2_1 U15033 ( .A(n11005), .B(n11023), .Y(n15590) );
  nand2_1 U15034 ( .A(n15792), .B(n15840), .Y(n11023) );
  and3_1 U15035 ( .A(n15715), .B(n15744), .C(n15714), .X(n15840) );
  nand3_1 U15036 ( .A(n15748), .B(n15833), .C(n15763), .Y(n11005) );
  inv_1 U15037 ( .A(n14302), .Y(n11009) );
  nor4_1 U15038 ( .A(n15842), .B(n15796), .C(n15680), .D(n15589), .Y(n15818)
         );
  nand2_1 U15039 ( .A(n14727), .B(n11024), .Y(n15589) );
  nand2_1 U15040 ( .A(n15778), .B(n15843), .Y(n11024) );
  nand3_1 U15041 ( .A(n15834), .B(n15786), .C(n15788), .Y(n14727) );
  inv_1 U15042 ( .A(n15844), .Y(n15786) );
  nand2_1 U15043 ( .A(n14762), .B(n14726), .Y(n15680) );
  nand2_1 U15044 ( .A(n15834), .B(n15843), .Y(n14726) );
  and3_1 U15045 ( .A(n15792), .B(n15779), .C(n15762), .X(n15843) );
  and2_0 U15046 ( .A(n15845), .B(n11314), .X(n15792) );
  and2_0 U15047 ( .A(n15806), .B(n15841), .X(n15834) );
  nand3_1 U15048 ( .A(n15778), .B(n15743), .C(n15765), .Y(n14762) );
  nor2_1 U15049 ( .A(n11319), .B(n15846), .Y(n15765) );
  nand4_1 U15050 ( .A(n14734), .B(n14737), .C(n14794), .D(n15847), .Y(n15796)
         );
  nor3_1 U15051 ( .A(n14825), .B(n15594), .C(n14782), .Y(n15847) );
  inv_1 U15052 ( .A(n14728), .Y(n14782) );
  nand2_1 U15053 ( .A(n15831), .B(n15752), .Y(n14728) );
  and2_0 U15054 ( .A(n15848), .B(n11314), .X(n15752) );
  and4_1 U15055 ( .A(n15829), .B(n15849), .C(n15743), .D(n24058), .X(n15831)
         );
  inv_1 U15056 ( .A(n10995), .Y(n15594) );
  nand2_1 U15057 ( .A(n15747), .B(n14780), .Y(n10995) );
  nand3_1 U15058 ( .A(n11030), .B(n15512), .C(n15551), .Y(n14825) );
  inv_1 U15059 ( .A(n15514), .Y(n15551) );
  nand2_1 U15060 ( .A(n14735), .B(n10989), .Y(n15514) );
  nand2_1 U15061 ( .A(n15850), .B(n15777), .Y(n10989) );
  nand2_1 U15062 ( .A(n14780), .B(n15777), .Y(n14735) );
  inv_1 U15063 ( .A(n15485), .Y(n14780) );
  nand4_1 U15064 ( .A(n15734), .B(n15719), .C(n15841), .D(n15743), .Y(n15512)
         );
  and2_0 U15065 ( .A(n15762), .B(n15851), .X(n15743) );
  nand3_1 U15066 ( .A(n15852), .B(n15777), .C(n15734), .Y(n11030) );
  nand3_1 U15067 ( .A(n15853), .B(n15718), .C(n15854), .Y(n14794) );
  nand3_1 U15068 ( .A(n15766), .B(n15753), .C(n15759), .Y(n14737) );
  and3_1 U15069 ( .A(n15754), .B(n15779), .C(n12916), .X(n15766) );
  nand2_1 U15070 ( .A(n15854), .B(n15761), .Y(n14734) );
  and3_1 U15071 ( .A(n15760), .B(n15798), .C(n15719), .X(n15854) );
  nand4_1 U15072 ( .A(n15780), .B(n14723), .C(n14738), .D(n15532), .Y(n15842)
         );
  nand2_1 U15073 ( .A(n15855), .B(n15742), .Y(n15532) );
  nand2_1 U15074 ( .A(n15855), .B(n15738), .Y(n14738) );
  and2_0 U15075 ( .A(n15856), .B(n15848), .X(n15738) );
  and3_1 U15076 ( .A(n15734), .B(n15829), .C(n15788), .X(n15855) );
  and2_0 U15077 ( .A(n15851), .B(n15798), .X(n15788) );
  inv_1 U15078 ( .A(n15857), .Y(n15829) );
  nand3_1 U15079 ( .A(n15776), .B(n15833), .C(n15744), .Y(n14723) );
  and2_0 U15080 ( .A(n15777), .B(n15745), .X(n15833) );
  nor2_1 U15081 ( .A(n15858), .B(n11442), .Y(n15777) );
  nor2_1 U15082 ( .A(n15846), .B(n11441), .Y(n15776) );
  nand3_1 U15083 ( .A(n15773), .B(n15745), .C(n15748), .Y(n15780) );
  nor2_1 U15084 ( .A(n11133), .B(n15718), .Y(n15748) );
  nor3_1 U15085 ( .A(n15859), .B(n15846), .C(n15860), .Y(n15773) );
  nand2_1 U15086 ( .A(inData[24]), .B(n14302), .Y(n10977) );
  nand3_1 U15087 ( .A(n14611), .B(n14636), .C(n14606), .Y(n14302) );
  and3_1 U15088 ( .A(n14708), .B(n14691), .C(n12472), .X(n14606) );
  inv_1 U15089 ( .A(n12355), .Y(n14691) );
  nor2_1 U15090 ( .A(n12316), .B(n24042), .Y(n14708) );
  nor2_1 U15091 ( .A(n14673), .B(n24045), .Y(n14636) );
  nor2_1 U15092 ( .A(n14701), .B(n14707), .Y(n14611) );
  and4_1 U15093 ( .A(n15861), .B(n15686), .C(n11001), .D(n15675), .X(n15817)
         );
  and4_1 U15094 ( .A(n14834), .B(n14763), .C(n15537), .D(n11003), .X(n15675)
         );
  nand4_1 U15095 ( .A(n15862), .B(n12916), .C(n12552), .D(n15863), .Y(n11003)
         );
  nand3_1 U15096 ( .A(n15751), .B(n15797), .C(n15862), .Y(n15537) );
  nor3_1 U15097 ( .A(n11400), .B(n15864), .C(n15865), .Y(n15862) );
  nand4_1 U15098 ( .A(n15717), .B(n15797), .C(n15751), .D(n15866), .Y(n14763)
         );
  nor2_1 U15099 ( .A(n15844), .B(n11400), .Y(n15866) );
  nand2_1 U15100 ( .A(n15867), .B(n15845), .Y(n15844) );
  inv_1 U15101 ( .A(n11500), .Y(n15797) );
  nand2_1 U15102 ( .A(n15816), .B(n15822), .Y(n14834) );
  and3_1 U15103 ( .A(n15764), .B(n15717), .C(n15755), .X(n15822) );
  and2_0 U15104 ( .A(n15798), .B(n15779), .X(n15755) );
  nor2_1 U15105 ( .A(n15718), .B(n11500), .Y(n15764) );
  inv_1 U15106 ( .A(n15864), .Y(n15816) );
  nand2_1 U15107 ( .A(n15856), .B(n15836), .Y(n15864) );
  nor2_1 U15108 ( .A(n15469), .B(n15784), .Y(n11001) );
  inv_1 U15109 ( .A(n15650), .Y(n15784) );
  nand3_1 U15110 ( .A(n15761), .B(n15717), .C(n15803), .Y(n15650) );
  nor2_1 U15111 ( .A(n15868), .B(n15718), .Y(n15761) );
  inv_1 U15112 ( .A(n14807), .Y(n15469) );
  nand4_1 U15113 ( .A(n15803), .B(n15853), .C(n15717), .D(n15718), .Y(n14807)
         );
  inv_1 U15114 ( .A(n15827), .Y(n15717) );
  and3_1 U15115 ( .A(n15815), .B(n15798), .C(n15763), .X(n15803) );
  and2_0 U15116 ( .A(n15867), .B(n15836), .X(n15763) );
  and4_1 U15117 ( .A(n10994), .B(n10992), .C(n14833), .D(n10991), .X(n15686)
         );
  nand4_1 U15118 ( .A(n15757), .B(n15789), .C(n15742), .D(n15744), .Y(n10991)
         );
  nor3_1 U15119 ( .A(n15795), .B(n24052), .C(n15718), .Y(n15744) );
  nor2_1 U15120 ( .A(n15869), .B(n15859), .Y(n15757) );
  nand4_1 U15121 ( .A(n15739), .B(n15735), .C(n15742), .D(n15745), .Y(n14833)
         );
  inv_1 U15122 ( .A(n15741), .Y(n15742) );
  nand2_1 U15123 ( .A(n15848), .B(n15867), .Y(n15741) );
  and2_0 U15124 ( .A(n15762), .B(n15870), .X(n15735) );
  nor2_1 U15125 ( .A(n15871), .B(n11444), .Y(n15762) );
  nand2_1 U15126 ( .A(n15458), .B(n15753), .Y(n10992) );
  nor3_1 U15127 ( .A(n10922), .B(n24055), .C(n15718), .Y(n15753) );
  and3_1 U15128 ( .A(n12916), .B(n15760), .C(n15712), .X(n15458) );
  and2_0 U15129 ( .A(n15835), .B(n15848), .X(n15712) );
  nor2_1 U15130 ( .A(n11445), .B(n24056), .Y(n15848) );
  nor2_1 U15131 ( .A(n15865), .B(n11211), .Y(n15760) );
  inv_1 U15132 ( .A(n15869), .Y(n12916) );
  nand4_1 U15133 ( .A(n15872), .B(n15759), .C(n15873), .D(n15789), .Y(n10994)
         );
  nor2_1 U15134 ( .A(n11500), .B(n15869), .Y(n15873) );
  inv_1 U15135 ( .A(n15812), .Y(n15759) );
  nand2_1 U15136 ( .A(n15835), .B(n15845), .Y(n15812) );
  and4_1 U15137 ( .A(n14817), .B(n15519), .C(n14791), .D(n15494), .X(n15861)
         );
  nand3_1 U15138 ( .A(n15789), .B(n15733), .C(n15807), .Y(n15494) );
  nor3_1 U15139 ( .A(n15868), .B(n11442), .C(n11400), .Y(n15807) );
  and2_0 U15140 ( .A(n15856), .B(n15845), .X(n15733) );
  nor2_1 U15141 ( .A(n11445), .B(n10613), .Y(n15845) );
  nand2_1 U15142 ( .A(n15850), .B(n14781), .Y(n14791) );
  inv_1 U15143 ( .A(n15484), .Y(n14781) );
  and3_1 U15144 ( .A(n15849), .B(n24058), .C(n15852), .X(n15850) );
  nand4_1 U15145 ( .A(n15789), .B(n15719), .C(n15739), .D(n15715), .Y(n15519)
         );
  nor2_1 U15146 ( .A(n15859), .B(n11442), .Y(n15715) );
  nor3_1 U15147 ( .A(n10832), .B(n24055), .C(n15718), .Y(n15739) );
  nor2_1 U15148 ( .A(n11320), .B(n15846), .Y(n15719) );
  inv_1 U15149 ( .A(n15615), .Y(n14817) );
  o21ai_0 U15150 ( .A1(n15484), .A2(n15485), .B1(n15495), .Y(n15615) );
  nand3_1 U15151 ( .A(n15734), .B(n15852), .C(n15747), .Y(n15495) );
  nor2_1 U15152 ( .A(n15869), .B(n15858), .Y(n15747) );
  nand2_1 U15153 ( .A(n24057), .B(n11444), .Y(n15869) );
  nor3_1 U15154 ( .A(n15857), .B(n15846), .C(n11443), .Y(n15852) );
  nand2_1 U15155 ( .A(n10613), .B(n11445), .Y(n15846) );
  nand4_1 U15156 ( .A(n24055), .B(n15718), .C(n12551), .D(n12550), .Y(n15857)
         );
  and2_0 U15157 ( .A(n15849), .B(n15874), .X(n15734) );
  nand3_1 U15158 ( .A(n15778), .B(n15836), .C(n15835), .Y(n15485) );
  nor2_1 U15159 ( .A(n10613), .B(n24059), .Y(n15836) );
  and3_1 U15160 ( .A(n15841), .B(n24058), .C(n15849), .X(n15778) );
  nor4_1 U15161 ( .A(n12550), .B(n12551), .C(n24051), .D(n24055), .Y(n15841)
         );
  nand2_1 U15162 ( .A(n15751), .B(n15779), .Y(n15484) );
  nor2_1 U15163 ( .A(n15875), .B(n24048), .Y(n15779) );
  nand2_1 U15164 ( .A(n15876), .B(n15877), .Y(n10350) );
  mux2i_1 U15165 ( .A0(n11847), .A1(n12506), .S(n11482), .Y(n15876) );
  inv_1 U15166 ( .A(n12564), .Y(n11847) );
  o32ai_1 U15167 ( .A1(n15878), .A2(n10609), .A3(n11086), .B1(n15879), .B2(
        n11775), .Y(n10349) );
  inv_1 U15168 ( .A(inData[14]), .Y(n11086) );
  o32ai_1 U15169 ( .A1(n15878), .A2(n15880), .A3(n11775), .B1(n15879), .B2(
        n15448), .Y(n10348) );
  inv_1 U15170 ( .A(inData[1]), .Y(n15448) );
  nand2_1 U15171 ( .A(n15881), .B(n10781), .Y(n10347) );
  nand2_1 U15172 ( .A(n15882), .B(n15879), .Y(n10781) );
  mux2i_1 U15173 ( .A0(n15883), .A1(n12826), .S(n10784), .Y(n15881) );
  xor2_1 U15174 ( .A(n15884), .B(n12331), .X(n15883) );
  o21ai_0 U15175 ( .A1(n15885), .A2(n15878), .B1(n15886), .Y(n10346) );
  nand2_1 U15176 ( .A(inData[3]), .B(n10784), .Y(n15886) );
  or2_0 U15177 ( .A(n15882), .B(n10784), .X(n15878) );
  inv_1 U15178 ( .A(n15879), .Y(n10784) );
  o211ai_1 U15179 ( .A1(n15887), .A2(n15888), .B1(n15889), .C1(n15890), .Y(
        n15879) );
  nor3_1 U15180 ( .A(n15891), .B(n23892), .C(n15892), .Y(n15882) );
  a21oi_1 U15181 ( .A1(n15893), .A2(n12331), .B1(n15894), .Y(n15885) );
  a21oi_1 U15182 ( .A1(n12331), .A2(n12408), .B1(n15895), .Y(n15894) );
  inv_1 U15183 ( .A(n15884), .Y(n15893) );
  nand2_1 U15184 ( .A(n15896), .B(n15897), .Y(n10345) );
  mux2i_1 U15185 ( .A0(n23958), .A1(n15898), .S(n15899), .Y(n15896) );
  nand2_1 U15186 ( .A(n15900), .B(n15897), .Y(n10344) );
  mux2i_1 U15187 ( .A0(n15901), .A1(n13958), .S(n15899), .Y(n15900) );
  inv_1 U15188 ( .A(inData[17]), .Y(n13958) );
  nand2_1 U15189 ( .A(inData[4]), .B(n15902), .Y(n15901) );
  o22ai_1 U15190 ( .A1(n10923), .A2(n15903), .B1(n15904), .B2(n15905), .Y(
        n10343) );
  xor2_1 U15191 ( .A(n1965), .B(n12393), .X(n15905) );
  nand2_1 U15192 ( .A(n15906), .B(n15897), .Y(n10342) );
  or2_0 U15193 ( .A(n15907), .B(n15899), .X(n15897) );
  mux2_1 U15194 ( .A0(n15908), .A1(inData[19]), .S(n15899), .X(n15906) );
  inv_1 U15195 ( .A(n15903), .Y(n15899) );
  xor2_1 U15196 ( .A(n15909), .B(n15910), .X(n15908) );
  mux2i_1 U15197 ( .A0(n15911), .A1(inData[4]), .S(n15912), .Y(n10341) );
  a211oi_1 U15198 ( .A1(n10608), .A2(n15913), .B1(n15914), .C1(n15915), .Y(
        n15911) );
  inv_1 U15199 ( .A(n15916), .Y(n15915) );
  o32ai_1 U15200 ( .A1(n15917), .A2(n10831), .A3(n15918), .B1(n12303), .B2(
        n15919), .Y(n10340) );
  inv_1 U15201 ( .A(inData[7]), .Y(n12303) );
  xor2_1 U15202 ( .A(n15920), .B(n15916), .X(n15917) );
  o22ai_1 U15203 ( .A1(n11355), .A2(n15919), .B1(n15921), .B2(n15918), .Y(
        n10339) );
  xor2_1 U15204 ( .A(n15916), .B(n23993), .X(n15921) );
  nor2_1 U15205 ( .A(n10774), .B(n10608), .Y(n10338) );
  o21ai_0 U15206 ( .A1(n10608), .A2(n15918), .B1(n15922), .Y(n10337) );
  nand2_1 U15207 ( .A(inData[5]), .B(n15912), .Y(n15922) );
  nand2_1 U15208 ( .A(n15923), .B(n15924), .Y(n10336) );
  mux2i_1 U15209 ( .A0(n15449), .A1(n15925), .S(n15926), .Y(n15923) );
  nand2_1 U15210 ( .A(inData[24]), .B(n15927), .Y(n15925) );
  xor2_1 U15211 ( .A(n15928), .B(n15929), .X(n15927) );
  nand2_1 U15212 ( .A(n12319), .B(n12302), .Y(n15929) );
  inv_1 U15213 ( .A(inData[23]), .Y(n15449) );
  o22ai_1 U15214 ( .A1(n15926), .A2(n12505), .B1(n23948), .B2(n15930), .Y(
        n10335) );
  o22ai_1 U15215 ( .A1(n14677), .A2(n15903), .B1(n15931), .B2(n15904), .Y(
        n10334) );
  inv_1 U15216 ( .A(inData[21]), .Y(n14677) );
  o32ai_1 U15217 ( .A1(n15904), .A2(n15932), .A3(n11367), .B1(n10831), .B2(
        n15903), .Y(n10333) );
  xor2_1 U15218 ( .A(n15933), .B(n12319), .X(n15932) );
  nand2_1 U15219 ( .A(n15907), .B(n15903), .Y(n15904) );
  o211ai_1 U15220 ( .A1(n15934), .A2(n15935), .B1(n15936), .C1(n15937), .Y(
        n15903) );
  a21oi_1 U15221 ( .A1(n15938), .A2(n15939), .B1(n15940), .Y(n15937) );
  nand3_1 U15222 ( .A(n15941), .B(n15934), .C(n15942), .Y(n15907) );
  a21oi_1 U15223 ( .A1(n15943), .A2(n23895), .B1(n15938), .Y(n15942) );
  nand2_1 U15224 ( .A(n15944), .B(n15924), .Y(n10332) );
  mux2_1 U15225 ( .A0(inData[25]), .A1(n15945), .S(n15926), .X(n15944) );
  nor2_1 U15226 ( .A(n23951), .B(n10831), .Y(n15945) );
  o32ai_1 U15227 ( .A1(n15898), .A2(n15946), .A3(n15930), .B1(n15926), .B2(
        n13959), .Y(n10331) );
  inv_1 U15228 ( .A(inData[27]), .Y(n13959) );
  xor2_1 U15229 ( .A(n15947), .B(n15948), .X(n15946) );
  nor2_1 U15230 ( .A(n12299), .B(n23951), .Y(n15948) );
  nand2_1 U15231 ( .A(n15949), .B(n15924), .Y(n10330) );
  nand4_1 U15232 ( .A(n15950), .B(n15926), .C(n15951), .D(n15952), .Y(n15924)
         );
  mux2i_1 U15233 ( .A0(n11545), .A1(n15953), .S(n15926), .Y(n15949) );
  o22ai_1 U15234 ( .A1(n15926), .A2(n12699), .B1(n15930), .B2(n15954), .Y(
        n10329) );
  xor2_1 U15235 ( .A(n15955), .B(n15956), .X(n15954) );
  nand2_1 U15236 ( .A(n15926), .B(n15957), .Y(n15930) );
  nand3_1 U15237 ( .A(n15951), .B(n15952), .C(n15950), .Y(n15957) );
  a211oi_1 U15238 ( .A1(n15184), .A2(n15958), .B1(n15959), .C1(n15960), .Y(
        n15926) );
  inv_1 U15239 ( .A(n15961), .Y(n15960) );
  a221oi_1 U15240 ( .A1(n15962), .A2(n15457), .B1(n15963), .B2(n15964), .C1(
        n15965), .Y(n15961) );
  nand2_1 U15241 ( .A(n15966), .B(n15967), .Y(n15964) );
  mux2i_1 U15242 ( .A0(n15967), .A1(n14873), .S(n23894), .Y(n15962) );
  o32ai_1 U15243 ( .A1(n15968), .A2(n23985), .A3(n15898), .B1(n11107), .B2(
        n15969), .Y(n10328) );
  o32ai_1 U15244 ( .A1(n15918), .A2(n15970), .A3(n11367), .B1(n12389), .B2(
        n15919), .Y(n10327) );
  inv_1 U15245 ( .A(inData[9]), .Y(n12389) );
  inv_1 U15246 ( .A(inData[8]), .Y(n11367) );
  nand2_1 U15247 ( .A(n15919), .B(n15971), .Y(n15918) );
  nor2_1 U15248 ( .A(n10774), .B(n15972), .Y(n10326) );
  nor2_1 U15249 ( .A(n10774), .B(n15970), .Y(n10325) );
  mux2i_1 U15250 ( .A0(n15973), .A1(inData[8]), .S(n15912), .Y(n10324) );
  inv_1 U15251 ( .A(n15919), .Y(n15912) );
  nand4_1 U15252 ( .A(n15974), .B(n15975), .C(n15976), .D(n15941), .Y(n15919)
         );
  o21ai_0 U15253 ( .A1(n15977), .A2(n15304), .B1(n15978), .Y(n15976) );
  mux2i_1 U15254 ( .A0(n15938), .A1(n15940), .S(n15939), .Y(n15974) );
  nor3_1 U15255 ( .A(n10831), .B(n15914), .C(n15979), .Y(n15973) );
  xor2_1 U15256 ( .A(n15972), .B(n15980), .X(n15979) );
  nor2_1 U15257 ( .A(n12401), .B(n15970), .Y(n15980) );
  inv_1 U15258 ( .A(n15971), .Y(n15914) );
  o211ai_1 U15259 ( .A1(n14873), .A2(n15981), .B1(n15982), .C1(n15983), .Y(
        n15971) );
  nor2_1 U15260 ( .A(n12401), .B(n10774), .Y(n10323) );
  mux2i_1 U15261 ( .A0(inData[11]), .A1(n15984), .S(n15969), .Y(n10322) );
  nor3_1 U15262 ( .A(n15985), .B(n15986), .C(n15898), .Y(n15984) );
  xor2_1 U15263 ( .A(n15987), .B(n15988), .X(n15985) );
  nor2_1 U15264 ( .A(n15972), .B(n15970), .Y(n15987) );
  mux2i_1 U15265 ( .A0(inData[14]), .A1(n15989), .S(n15969), .Y(n10321) );
  nor2_1 U15266 ( .A(n15986), .B(n15990), .Y(n15989) );
  inv_1 U15267 ( .A(n15991), .Y(n15986) );
  o32ai_1 U15268 ( .A1(n15968), .A2(n23981), .A3(n12699), .B1(n13374), .B2(
        n15969), .Y(n10320) );
  inv_1 U15269 ( .A(inData[13]), .Y(n13374) );
  nor2_1 U15270 ( .A(n15992), .B(n12628), .Y(n10319) );
  o22ai_1 U15271 ( .A1(n15969), .A2(n15993), .B1(n15994), .B2(n15968), .Y(
        n10318) );
  xor2_1 U15272 ( .A(n15992), .B(n15995), .X(n15994) );
  o32ai_1 U15273 ( .A1(n15968), .A2(n15996), .A3(n11134), .B1(n15969), .B2(
        n15997), .Y(n10317) );
  inv_1 U15274 ( .A(inData[15]), .Y(n15997) );
  a21oi_1 U15275 ( .A1(n15995), .A2(n12394), .B1(n15998), .Y(n15996) );
  a21oi_1 U15276 ( .A1(n12394), .A2(n15999), .B1(n16000), .Y(n15998) );
  inv_1 U15277 ( .A(n16001), .Y(n15995) );
  nand2_1 U15278 ( .A(n15969), .B(n15991), .Y(n15968) );
  nand3_1 U15279 ( .A(n15983), .B(n15936), .C(n15950), .Y(n15991) );
  nand4_1 U15280 ( .A(n15936), .B(n15952), .C(n16002), .D(n16003), .Y(n15969)
         );
  a221oi_1 U15281 ( .A1(n16004), .A2(n23893), .B1(n15978), .B2(n23894), .C1(
        n15940), .Y(n16003) );
  nand2_1 U15282 ( .A(n15887), .B(n16005), .Y(n15940) );
  nand2_1 U15283 ( .A(n12636), .B(n15999), .Y(n10316) );
  o32ai_1 U15284 ( .A1(n16006), .A2(n16007), .A3(n12826), .B1(n16008), .B2(
        n11134), .Y(n10315) );
  mux2i_1 U15285 ( .A0(inData[29]), .A1(n16009), .S(n16008), .Y(n10314) );
  and3_1 U15286 ( .A(inData[4]), .B(n16010), .C(n23949), .X(n16009) );
  o32ai_1 U15287 ( .A1(n16011), .A2(n11330), .A3(n16006), .B1(n16008), .B2(
        n11175), .Y(n10313) );
  xor2_1 U15288 ( .A(n23950), .B(n23949), .X(n16011) );
  o32ai_1 U15289 ( .A1(n16006), .A2(n16012), .A3(n11107), .B1(n16008), .B2(
        n13954), .Y(n10312) );
  inv_1 U15290 ( .A(inData[31]), .Y(n13954) );
  xor2_1 U15291 ( .A(n16013), .B(n16014), .X(n16012) );
  nor2_1 U15292 ( .A(n23950), .B(n16015), .Y(n16014) );
  nand2_1 U15293 ( .A(n16008), .B(n16010), .Y(n16006) );
  o21ai_0 U15294 ( .A1(n23871), .A2(n24036), .B1(n15362), .Y(n16010) );
  inv_1 U15295 ( .A(n23873), .Y(n15362) );
  and2_0 U15296 ( .A(n16016), .B(n16017), .X(n16008) );
  o21ai_0 U15297 ( .A1(n23873), .A2(n15398), .B1(n23872), .Y(n16017) );
  inv_1 U15298 ( .A(n23871), .Y(n15398) );
  xor2_1 U15299 ( .A(n16018), .B(n23873), .X(n16016) );
  nand2_1 U15300 ( .A(n23871), .B(n24036), .Y(n16018) );
  o21ai_0 U15301 ( .A1(n16019), .A2(n10683), .B1(n16020), .Y(n10311) );
  mux2i_1 U15302 ( .A0(n10685), .A1(n16021), .S(n16022), .Y(n16020) );
  nor4_1 U15303 ( .A(n16023), .B(n14266), .C(n14055), .D(n14148), .Y(n16022)
         );
  nand4_1 U15304 ( .A(n14046), .B(n10696), .C(n14007), .D(n16024), .Y(n14148)
         );
  and3_1 U15305 ( .A(n13969), .B(n14040), .C(n14177), .X(n16024) );
  inv_1 U15306 ( .A(n14172), .Y(n14055) );
  nand3_1 U15307 ( .A(n16025), .B(n14139), .C(n16026), .Y(n14266) );
  and3_1 U15308 ( .A(n12774), .B(n10710), .C(n10700), .X(n16026) );
  inv_1 U15309 ( .A(n16027), .Y(n16025) );
  nand4_1 U15310 ( .A(n14157), .B(n12777), .C(n14153), .D(n14057), .Y(n16023)
         );
  nor4_1 U15311 ( .A(n16028), .B(n16029), .C(n14130), .D(n16030), .Y(n16021)
         );
  nand3_1 U15312 ( .A(n14018), .B(n10727), .C(n14033), .Y(n14130) );
  nand3_1 U15313 ( .A(n12773), .B(n14143), .C(n14205), .Y(n16029) );
  inv_1 U15314 ( .A(n10705), .Y(n14205) );
  nand2_1 U15315 ( .A(n14187), .B(n14218), .Y(n10705) );
  nand4_1 U15316 ( .A(n16031), .B(n16032), .C(n16033), .D(n16034), .Y(n14143)
         );
  and4_1 U15317 ( .A(n10727), .B(n14245), .C(n14219), .D(n14033), .X(n16034)
         );
  nand2_1 U15318 ( .A(n16035), .B(n16036), .Y(n14033) );
  nand3_1 U15319 ( .A(n16037), .B(n16038), .C(n16039), .Y(n14219) );
  nand3_1 U15320 ( .A(n16040), .B(n16041), .C(n16042), .Y(n10727) );
  nor4_1 U15321 ( .A(n14147), .B(n10690), .C(n16027), .D(n14223), .Y(n16033)
         );
  nand3_1 U15322 ( .A(n16043), .B(n14188), .C(n16044), .Y(n14223) );
  and4_1 U15323 ( .A(n13978), .B(n14172), .C(n14017), .D(n13985), .X(n16044)
         );
  nand4_1 U15324 ( .A(n16045), .B(n16046), .C(n16047), .D(n16048), .Y(n13985)
         );
  nand4_1 U15325 ( .A(n16049), .B(n16050), .C(n16046), .D(n16051), .Y(n14017)
         );
  nand4_1 U15326 ( .A(n16040), .B(n16052), .C(n23962), .D(n16053), .Y(n14172)
         );
  nand3_1 U15327 ( .A(n16054), .B(n16055), .C(n16056), .Y(n13978) );
  and4_1 U15328 ( .A(n14052), .B(n13974), .C(n10725), .D(n16057), .X(n14188)
         );
  nand3_1 U15329 ( .A(n16058), .B(n16059), .C(n16060), .Y(n10725) );
  nand3_1 U15330 ( .A(n16058), .B(n16061), .C(n16042), .Y(n13974) );
  nand3_1 U15331 ( .A(n16039), .B(n16062), .C(n16049), .Y(n14052) );
  a21oi_1 U15332 ( .A1(n16063), .A2(n16064), .B1(n14082), .Y(n16043) );
  nand4_1 U15333 ( .A(n12772), .B(n14050), .C(n14177), .D(n10694), .Y(n14082)
         );
  nand2_1 U15334 ( .A(n16065), .B(n16066), .Y(n10694) );
  nand3_1 U15335 ( .A(n16067), .B(n16068), .C(n16069), .Y(n14177) );
  nand3_1 U15336 ( .A(n16070), .B(n16071), .C(n16067), .Y(n14050) );
  nand3_1 U15337 ( .A(n16038), .B(n16054), .C(n16061), .Y(n12772) );
  nand3_1 U15338 ( .A(n13976), .B(n12759), .C(n14114), .Y(n16027) );
  nor2_1 U15339 ( .A(n12752), .B(n12844), .Y(n14114) );
  inv_1 U15340 ( .A(n10697), .Y(n12844) );
  nand2_1 U15341 ( .A(n16055), .B(n16036), .Y(n10697) );
  nand2_1 U15342 ( .A(n10695), .B(n14060), .Y(n12752) );
  nand2_1 U15343 ( .A(n16072), .B(n16073), .Y(n14060) );
  nand3_1 U15344 ( .A(n16074), .B(n16075), .C(n16076), .Y(n10695) );
  nand3_1 U15345 ( .A(n16077), .B(n16058), .C(n16037), .Y(n12759) );
  nand3_1 U15346 ( .A(n16042), .B(n16077), .C(n16078), .Y(n13976) );
  nand4_1 U15347 ( .A(n13979), .B(n14024), .C(n16079), .D(n16080), .Y(n10690)
         );
  and4_1 U15348 ( .A(n14093), .B(n14062), .C(n14139), .D(n13969), .X(n16080)
         );
  inv_1 U15349 ( .A(n16081), .Y(n13969) );
  o21ai_0 U15350 ( .A1(n14215), .A2(n14216), .B1(n14267), .Y(n16081) );
  nand3_1 U15351 ( .A(n16082), .B(n16075), .C(n16061), .Y(n14267) );
  and2_0 U15352 ( .A(n16083), .B(n16071), .X(n16061) );
  and3_1 U15353 ( .A(n12775), .B(n14180), .C(n14221), .X(n14139) );
  nand4_1 U15354 ( .A(n16037), .B(n16050), .C(n16058), .D(n16084), .Y(n14221)
         );
  nand3_1 U15355 ( .A(n16056), .B(n16046), .C(n16041), .Y(n14180) );
  nand3_1 U15356 ( .A(n16067), .B(n16066), .C(n16069), .Y(n12775) );
  nand4_1 U15357 ( .A(n16085), .B(n16086), .C(n16087), .D(n16088), .Y(n14062)
         );
  nand3_1 U15358 ( .A(n16086), .B(n16089), .C(n16090), .Y(n14093) );
  and3_1 U15359 ( .A(n12777), .B(n14046), .C(n14153), .X(n16079) );
  nand3_1 U15360 ( .A(n16091), .B(n16055), .C(n16090), .Y(n14153) );
  nand4_1 U15361 ( .A(n16046), .B(n16068), .C(n16092), .D(n16093), .Y(n14046)
         );
  nand2_1 U15362 ( .A(n16058), .B(n16094), .Y(n12777) );
  nand4_1 U15363 ( .A(n16035), .B(n16095), .C(n16087), .D(n16088), .Y(n14024)
         );
  nand3_1 U15364 ( .A(n16046), .B(n16047), .C(n16077), .Y(n13979) );
  inv_1 U15365 ( .A(n12760), .Y(n14147) );
  nand2_1 U15366 ( .A(n16096), .B(n16063), .Y(n12760) );
  nor4_1 U15367 ( .A(n14248), .B(n14242), .C(n12753), .D(n14225), .Y(n16032)
         );
  nand4_1 U15368 ( .A(n14081), .B(n12778), .C(n16097), .D(n16098), .Y(n14225)
         );
  and4_1 U15369 ( .A(n14065), .B(n14051), .C(n14018), .D(n14016), .X(n16098)
         );
  nor3_1 U15370 ( .A(n14270), .B(n10715), .C(n14262), .Y(n14016) );
  inv_1 U15371 ( .A(n14098), .Y(n14262) );
  inv_1 U15372 ( .A(n14077), .Y(n10715) );
  inv_1 U15373 ( .A(n10719), .Y(n14270) );
  nand4_1 U15374 ( .A(n16099), .B(n16100), .C(n16101), .D(n16102), .Y(n10719)
         );
  nor2_1 U15375 ( .A(n16103), .B(n16104), .Y(n16102) );
  nand3_1 U15376 ( .A(n16105), .B(n16047), .C(n16069), .Y(n14018) );
  nand3_1 U15377 ( .A(n16056), .B(n16035), .C(n16037), .Y(n14051) );
  nand4_1 U15378 ( .A(n16106), .B(n16099), .C(n16107), .D(n16108), .Y(n14065)
         );
  and2_0 U15379 ( .A(n16062), .B(n16068), .X(n16108) );
  and2_0 U15380 ( .A(n14104), .B(n14029), .X(n16097) );
  nand3_1 U15381 ( .A(n16067), .B(n16095), .C(n16049), .Y(n12778) );
  nand4_1 U15382 ( .A(n14115), .B(n14204), .C(n12771), .D(n16109), .Y(n12753)
         );
  and4_1 U15383 ( .A(n10718), .B(n10720), .C(n14006), .D(n14080), .X(n16109)
         );
  nand4_1 U15384 ( .A(n16078), .B(n16073), .C(n16084), .D(n16110), .Y(n14080)
         );
  nand3_1 U15385 ( .A(n16111), .B(n16112), .C(n16058), .Y(n14006) );
  inv_1 U15386 ( .A(n16104), .Y(n16058) );
  nand2_1 U15387 ( .A(n16113), .B(n23962), .Y(n16104) );
  nand3_1 U15388 ( .A(n16111), .B(n16051), .C(n16038), .Y(n10718) );
  and2_0 U15389 ( .A(n13975), .B(n14001), .X(n14204) );
  nand2_1 U15390 ( .A(n16114), .B(n16066), .Y(n14001) );
  and3_1 U15391 ( .A(n14227), .B(n14179), .C(n16115), .X(n14115) );
  and3_1 U15392 ( .A(n14005), .B(n14097), .C(n14218), .X(n16115) );
  nand3_1 U15393 ( .A(n16076), .B(n16116), .C(n16111), .Y(n14218) );
  nand4_1 U15394 ( .A(n16051), .B(n16086), .C(n16054), .D(n16110), .Y(n14097)
         );
  nand2_1 U15395 ( .A(n16117), .B(n16118), .Y(n14005) );
  and3_1 U15396 ( .A(n13999), .B(n10696), .C(n13968), .X(n14179) );
  inv_1 U15397 ( .A(n10691), .Y(n13968) );
  nand2_1 U15398 ( .A(n14057), .B(n14207), .Y(n10691) );
  nand3_1 U15399 ( .A(n16112), .B(n16118), .C(n16047), .Y(n14207) );
  nand2_1 U15400 ( .A(n16111), .B(n16117), .Y(n14057) );
  and4_1 U15401 ( .A(n16107), .B(n16119), .C(n16120), .D(n16116), .X(n16117)
         );
  nor2_1 U15402 ( .A(n23974), .B(n23962), .Y(n16120) );
  inv_1 U15403 ( .A(n16121), .Y(n16119) );
  nand2_1 U15404 ( .A(n16075), .B(n16122), .Y(n10696) );
  nand3_1 U15405 ( .A(n16118), .B(n16084), .C(n16049), .Y(n13999) );
  and2_0 U15406 ( .A(n16123), .B(n16100), .X(n16118) );
  and4_1 U15407 ( .A(n13988), .B(n14000), .C(n14007), .D(n10699), .X(n14227)
         );
  nand3_1 U15408 ( .A(n16111), .B(n16089), .C(n16035), .Y(n14007) );
  nand2_1 U15409 ( .A(n16078), .B(n16114), .Y(n14000) );
  nand4_1 U15410 ( .A(n16086), .B(n16124), .C(n16074), .D(n16075), .Y(n13988)
         );
  nand2_1 U15411 ( .A(n14157), .B(n10726), .Y(n14242) );
  nand2_1 U15412 ( .A(n16125), .B(n16055), .Y(n10726) );
  nand3_1 U15413 ( .A(n16126), .B(n16127), .C(n16052), .Y(n14157) );
  nand4_1 U15414 ( .A(n12774), .B(n14019), .C(n16128), .D(n16129), .Y(n14248)
         );
  nor4_1 U15415 ( .A(n13990), .B(n13995), .C(n16130), .D(n16131), .Y(n16129)
         );
  inv_1 U15416 ( .A(n14178), .Y(n13995) );
  nand3_1 U15417 ( .A(n16112), .B(n16059), .C(n16035), .Y(n14178) );
  and2_0 U15418 ( .A(n16107), .B(n16093), .X(n16112) );
  inv_1 U15419 ( .A(n14117), .Y(n13990) );
  nand3_1 U15420 ( .A(n16035), .B(n16075), .C(n16077), .Y(n14117) );
  and2_0 U15421 ( .A(n16051), .B(n16048), .X(n16077) );
  and3_1 U15422 ( .A(n10692), .B(n16132), .C(n10710), .X(n16128) );
  nand3_1 U15423 ( .A(n16041), .B(n16052), .C(n16133), .Y(n10710) );
  nand3_1 U15424 ( .A(n16070), .B(n16134), .C(n16062), .Y(n10692) );
  and3_1 U15425 ( .A(n16048), .B(n16116), .C(n16038), .X(n16070) );
  nand4_1 U15426 ( .A(n16050), .B(n16107), .C(n16135), .D(n16116), .Y(n12774)
         );
  nor3_1 U15427 ( .A(n12785), .B(n14201), .C(n10723), .Y(n16031) );
  nand4_1 U15428 ( .A(n14138), .B(n14003), .C(n14056), .D(n14092), .Y(n10723)
         );
  nand2_1 U15429 ( .A(n16125), .B(n16063), .Y(n14056) );
  inv_1 U15430 ( .A(n14165), .Y(n14138) );
  nand2_1 U15431 ( .A(n14090), .B(n16136), .Y(n14165) );
  nand4_1 U15432 ( .A(n16050), .B(n16071), .C(n16137), .D(n16138), .Y(n16136)
         );
  nor3_1 U15433 ( .A(n16139), .B(n16140), .C(n16141), .Y(n16138) );
  nand3_1 U15434 ( .A(n16067), .B(n16085), .C(n16063), .Y(n14090) );
  nand4_1 U15435 ( .A(n14040), .B(n14187), .C(n10700), .D(n10709), .Y(n12785)
         );
  nand2_1 U15436 ( .A(n16135), .B(n16126), .Y(n10700) );
  nand3_1 U15437 ( .A(n16090), .B(n16082), .C(n16060), .Y(n14187) );
  nand3_1 U15438 ( .A(n16047), .B(n16052), .C(n16069), .Y(n14040) );
  and2_0 U15439 ( .A(n16060), .B(n16048), .X(n16069) );
  inv_1 U15440 ( .A(n14169), .Y(n12773) );
  nand2_1 U15441 ( .A(n14245), .B(n16132), .Y(n14169) );
  nand4_1 U15442 ( .A(n16041), .B(n16090), .C(n16107), .D(n16106), .Y(n16132)
         );
  nand3_1 U15443 ( .A(n16133), .B(n16105), .C(n16063), .Y(n14245) );
  nand4_1 U15444 ( .A(n14003), .B(n12757), .C(n10720), .D(n16142), .Y(n16028)
         );
  and2_0 U15445 ( .A(n14098), .B(n13975), .X(n16142) );
  nand4_1 U15446 ( .A(n16042), .B(n16035), .C(n16143), .D(n16110), .Y(n13975)
         );
  nand3_1 U15447 ( .A(n16035), .B(n16073), .C(n16085), .Y(n14098) );
  and2_0 U15448 ( .A(n16092), .B(n16106), .X(n16085) );
  nand4_1 U15449 ( .A(n16041), .B(n16084), .C(n16075), .D(n16110), .Y(n10720)
         );
  nor2_1 U15450 ( .A(n16140), .B(n16144), .Y(n16075) );
  nand2_1 U15451 ( .A(n16125), .B(n16035), .Y(n14003) );
  and2_0 U15452 ( .A(n16126), .B(n16145), .X(n16125) );
  and3_1 U15453 ( .A(n16048), .B(n16071), .C(n16106), .X(n16126) );
  inv_1 U15454 ( .A(n12750), .Y(n10685) );
  nand2_1 U15455 ( .A(inData[11]), .B(n12757), .Y(n12750) );
  inv_1 U15456 ( .A(n14164), .Y(n10683) );
  nor2_1 U15457 ( .A(n12747), .B(inData[11]), .Y(n14164) );
  inv_1 U15458 ( .A(n12757), .Y(n12747) );
  nand3_1 U15459 ( .A(n13831), .B(n13832), .C(n13837), .Y(n12757) );
  inv_1 U15460 ( .A(n16146), .Y(n13837) );
  nor2_1 U15461 ( .A(n16147), .B(n23903), .Y(n13832) );
  inv_1 U15462 ( .A(n16148), .Y(n13831) );
  inv_1 U15463 ( .A(n16030), .Y(n16019) );
  nand4_1 U15464 ( .A(n14104), .B(n14092), .C(n16149), .D(n16150), .Y(n16030)
         );
  nor4_1 U15465 ( .A(n14201), .B(n16151), .C(n14170), .D(n14069), .Y(n16150)
         );
  nand4_1 U15466 ( .A(n14081), .B(n14025), .C(n14029), .D(n16152), .Y(n14069)
         );
  nor2_1 U15467 ( .A(n16131), .B(n10722), .Y(n16152) );
  nand2_1 U15468 ( .A(n14019), .B(n16057), .Y(n10722) );
  nand3_1 U15469 ( .A(n16153), .B(n16055), .C(n16105), .Y(n16057) );
  nand3_1 U15470 ( .A(n16091), .B(n16059), .C(n16078), .Y(n14019) );
  nor2_1 U15471 ( .A(n16154), .B(n16155), .Y(n16078) );
  inv_1 U15472 ( .A(n16103), .Y(n16091) );
  nand4_1 U15473 ( .A(n12751), .B(n10717), .C(n14108), .D(n10707), .Y(n16131)
         );
  nand3_1 U15474 ( .A(n16050), .B(n16062), .C(n16156), .Y(n10707) );
  nor3_1 U15475 ( .A(n16157), .B(n16158), .C(n16159), .Y(n16156) );
  nand3_1 U15476 ( .A(n16056), .B(n16052), .C(n16063), .Y(n14108) );
  and2_0 U15477 ( .A(n16045), .B(n16099), .X(n16056) );
  nand3_1 U15478 ( .A(n16133), .B(n16067), .C(n16049), .Y(n10717) );
  inv_1 U15479 ( .A(n16160), .Y(n16133) );
  nand4_1 U15480 ( .A(n16050), .B(n16051), .C(n16161), .D(n16101), .Y(n12751)
         );
  and2_0 U15481 ( .A(n16162), .B(n16055), .X(n16161) );
  nand2_1 U15482 ( .A(n16096), .B(n16049), .Y(n14029) );
  nor3_1 U15483 ( .A(n16163), .B(n23962), .C(n16164), .Y(n16049) );
  and3_1 U15484 ( .A(n16143), .B(n16099), .C(n16037), .X(n16096) );
  nand2_1 U15485 ( .A(n16063), .B(n16064), .Y(n14025) );
  o32ai_1 U15486 ( .A1(n16165), .A2(n16166), .A3(n16103), .B1(n16167), .B2(
        n16160), .Y(n16064) );
  nand2_1 U15487 ( .A(n16093), .B(n16134), .Y(n16103) );
  nand2_1 U15488 ( .A(n16094), .B(n16066), .Y(n14081) );
  and3_1 U15489 ( .A(n16153), .B(n16168), .C(n16101), .X(n16094) );
  nand2_1 U15490 ( .A(n14061), .B(n14263), .Y(n14170) );
  nand4_1 U15491 ( .A(n16067), .B(n16050), .C(n16082), .D(n16084), .Y(n14263)
         );
  nand2_1 U15492 ( .A(n16065), .B(n16082), .Y(n14061) );
  nand2_1 U15493 ( .A(n16169), .B(n12771), .Y(n16151) );
  and4_1 U15494 ( .A(n14137), .B(n14116), .C(n14123), .D(n14078), .X(n12771)
         );
  nand4_1 U15495 ( .A(n16123), .B(n16162), .C(n16076), .D(n16116), .Y(n14078)
         );
  nand4_1 U15496 ( .A(n16042), .B(n16045), .C(n16038), .D(n16110), .Y(n14123)
         );
  nor2_1 U15497 ( .A(n16170), .B(n16144), .Y(n16042) );
  inv_1 U15498 ( .A(n14244), .Y(n14116) );
  nand2_1 U15499 ( .A(n13987), .B(n13996), .Y(n14244) );
  nand2_1 U15500 ( .A(n16054), .B(n16122), .Y(n13996) );
  and4_1 U15501 ( .A(n23962), .B(n16053), .C(n16110), .D(n16089), .X(n16122)
         );
  nor2_1 U15502 ( .A(n16141), .B(n16171), .Y(n16089) );
  nand3_1 U15503 ( .A(n16038), .B(n16111), .C(n16045), .Y(n13987) );
  and3_1 U15504 ( .A(n16172), .B(n16110), .C(n16087), .X(n16111) );
  and2_0 U15505 ( .A(n16173), .B(n16155), .X(n16038) );
  and2_0 U15506 ( .A(n10693), .B(n10706), .X(n14137) );
  nand2_1 U15507 ( .A(n16114), .B(n16041), .Y(n10706) );
  nor3_1 U15508 ( .A(n16163), .B(n16155), .C(n16164), .Y(n16041) );
  and4_1 U15509 ( .A(n16087), .B(n16172), .C(n16074), .D(n16071), .X(n16114)
         );
  nor3_1 U15510 ( .A(n16174), .B(n11520), .C(n16175), .Y(n16074) );
  nand4_1 U15511 ( .A(n16051), .B(n16123), .C(n16086), .D(n16162), .Y(n10693)
         );
  inv_1 U15512 ( .A(n16157), .Y(n16086) );
  nand2_1 U15513 ( .A(n16173), .B(n23962), .Y(n16157) );
  and2_0 U15514 ( .A(n16101), .B(n16110), .X(n16123) );
  nor2_1 U15515 ( .A(n16176), .B(n16177), .Y(n16051) );
  inv_1 U15516 ( .A(n16130), .Y(n16169) );
  nand4_1 U15517 ( .A(n14102), .B(n14171), .C(n10701), .D(n10708), .Y(n16130)
         );
  inv_1 U15518 ( .A(n14106), .Y(n10708) );
  nor2_1 U15519 ( .A(n16167), .B(n14216), .Y(n14106) );
  nand3_1 U15520 ( .A(n16048), .B(n16055), .C(n16045), .Y(n14216) );
  nor2_1 U15521 ( .A(n16178), .B(n23962), .Y(n16055) );
  nand3_1 U15522 ( .A(n16082), .B(n16153), .C(n16052), .Y(n10701) );
  nor2_1 U15523 ( .A(n16179), .B(n16180), .Y(n16052) );
  and2_0 U15524 ( .A(n16143), .B(n16048), .X(n16153) );
  and2_0 U15525 ( .A(n16113), .B(n16155), .X(n16082) );
  nand3_1 U15526 ( .A(n16095), .B(n16047), .C(n16067), .Y(n14171) );
  nor2_1 U15527 ( .A(n16179), .B(n16170), .Y(n16067) );
  nor2_1 U15528 ( .A(n16154), .B(n23962), .Y(n16047) );
  nor3_1 U15529 ( .A(n16176), .B(n16159), .C(n16165), .Y(n16095) );
  nand3_1 U15530 ( .A(n16059), .B(n16066), .C(n16060), .Y(n14102) );
  nor2_1 U15531 ( .A(n16175), .B(n16171), .Y(n16060) );
  nand4_1 U15532 ( .A(n14045), .B(n14004), .C(n14166), .D(n14101), .Y(n14201)
         );
  nand2_1 U15533 ( .A(n16063), .B(n16065), .Y(n14101) );
  nor2_1 U15534 ( .A(n16160), .B(n16166), .Y(n16065) );
  nand3_1 U15535 ( .A(n16106), .B(n16099), .C(n16124), .Y(n16160) );
  nand3_1 U15536 ( .A(n16063), .B(n16046), .C(n16039), .Y(n14166) );
  and2_0 U15537 ( .A(n16050), .B(n16143), .X(n16039) );
  nor2_1 U15538 ( .A(n16159), .B(n16171), .Y(n16143) );
  inv_1 U15539 ( .A(n16165), .Y(n16050) );
  nand2_1 U15540 ( .A(n16181), .B(n11520), .Y(n16165) );
  inv_1 U15541 ( .A(n16182), .Y(n16046) );
  nand4_1 U15542 ( .A(n16035), .B(n16105), .C(n16092), .D(n16183), .Y(n14004)
         );
  nor2_1 U15543 ( .A(n16139), .B(n23962), .Y(n16035) );
  nand3_1 U15544 ( .A(n16068), .B(n16062), .C(n16040), .Y(n14045) );
  and2_0 U15545 ( .A(n16083), .B(n16124), .X(n16040) );
  nor3_1 U15546 ( .A(n10615), .B(n12297), .C(n16184), .Y(n16083) );
  and3_1 U15547 ( .A(n14077), .B(n10709), .C(n10699), .X(n16149) );
  nand2_1 U15548 ( .A(n16054), .B(n16072), .Y(n10699) );
  and3_1 U15549 ( .A(n16076), .B(n16110), .C(n16106), .X(n16072) );
  inv_1 U15550 ( .A(n16159), .Y(n16106) );
  nor3_1 U15551 ( .A(n11520), .B(n24006), .C(n10615), .Y(n16110) );
  and2_0 U15552 ( .A(n16066), .B(n16071), .X(n16076) );
  nor3_1 U15553 ( .A(n16155), .B(n23974), .C(n16121), .Y(n16066) );
  inv_1 U15554 ( .A(n14215), .Y(n16054) );
  nand3_1 U15555 ( .A(n16068), .B(n16048), .C(n16185), .Y(n10709) );
  nor3_1 U15556 ( .A(n16186), .B(n16158), .C(n16175), .Y(n16185) );
  nor2_1 U15557 ( .A(n16178), .B(n16155), .Y(n16068) );
  nand2_1 U15558 ( .A(n16127), .B(n16036), .Y(n14077) );
  and2_0 U15559 ( .A(n16084), .B(n16059), .X(n16036) );
  and2_0 U15560 ( .A(n16145), .B(n16099), .X(n16059) );
  inv_1 U15561 ( .A(n16186), .Y(n16145) );
  nor2_1 U15562 ( .A(n16177), .B(n16158), .Y(n16084) );
  nand3_1 U15563 ( .A(n16135), .B(n16183), .C(n16092), .Y(n14092) );
  and2_0 U15564 ( .A(n16107), .B(n16048), .X(n16092) );
  nor2_1 U15565 ( .A(n16187), .B(n12297), .Y(n16048) );
  and2_0 U15566 ( .A(n16073), .B(n16127), .X(n16135) );
  nor2_1 U15567 ( .A(n16188), .B(n23962), .Y(n16127) );
  nor2_1 U15568 ( .A(n16189), .B(n16170), .Y(n16073) );
  nand3_1 U15569 ( .A(n16090), .B(n16045), .C(n16063), .Y(n14104) );
  nor2_1 U15570 ( .A(n16188), .B(n16155), .Y(n16063) );
  nor2_1 U15571 ( .A(n16176), .B(n16141), .Y(n16045) );
  and2_0 U15572 ( .A(n16105), .B(n16099), .X(n16090) );
  nor2_1 U15573 ( .A(n16190), .B(n12297), .Y(n16099) );
  inv_1 U15574 ( .A(n16191), .Y(n16105) );
  mux2i_1 U15575 ( .A0(n16192), .A1(n16193), .S(n12586), .Y(n10310) );
  nand2_1 U15576 ( .A(n23922), .B(n16194), .Y(n16193) );
  xor2_1 U15577 ( .A(n16195), .B(n16196), .X(n16194) );
  mux2i_1 U15578 ( .A0(n11567), .A1(n11566), .S(n16195), .Y(n16192) );
  nor2_1 U15579 ( .A(n10774), .B(n16197), .Y(n11566) );
  nor2_1 U15580 ( .A(n16198), .B(n10774), .Y(n11567) );
  nand2_1 U15581 ( .A(n23922), .B(n16199), .Y(n10309) );
  xnor2_1 U15582 ( .A(n34), .B(n16200), .Y(n16199) );
  nand2_1 U15583 ( .A(n16201), .B(n16202), .Y(n16200) );
  inv_1 U15584 ( .A(n16203), .Y(n16201) );
  mux2i_1 U15585 ( .A0(n16204), .A1(n16205), .S(n11152), .Y(n10308) );
  nand2_1 U15586 ( .A(n16206), .B(n11150), .Y(n11152) );
  nor3_1 U15587 ( .A(n11175), .B(n16207), .C(n11150), .Y(n16205) );
  xor2_1 U15588 ( .A(n16208), .B(n20750), .X(n16207) );
  nand2_1 U15589 ( .A(n23928), .B(n12376), .Y(n16208) );
  xor2_1 U15590 ( .A(n16209), .B(n16210), .X(n16204) );
  xor2_1 U15591 ( .A(n23909), .B(n16211), .X(n16210) );
  o21ai_0 U15592 ( .A1(n11213), .A2(n16212), .B1(n16213), .Y(n10307) );
  mux2i_1 U15593 ( .A0(n11267), .A1(n11266), .S(n63), .Y(n16213) );
  inv_1 U15594 ( .A(n11289), .Y(n11266) );
  o21ai_0 U15595 ( .A1(n11288), .A2(n11212), .B1(n15815), .Y(n11289) );
  nor3_1 U15596 ( .A(n11212), .B(n11288), .C(n11211), .Y(n11267) );
  xor2_1 U15597 ( .A(n16214), .B(n16215), .X(n16212) );
  xor2_1 U15598 ( .A(n10942), .B(n16216), .X(n16215) );
  xor2_1 U15599 ( .A(n5), .B(n16217), .X(n16214) );
  nor2_1 U15600 ( .A(n16218), .B(n10774), .Y(n10306) );
  xor2_1 U15601 ( .A(n10862), .B(n16219), .X(n16218) );
  xor2_1 U15602 ( .A(n23801), .B(n10813), .X(n16219) );
  mux2i_1 U15603 ( .A0(n16220), .A1(n16221), .S(n16222), .Y(n10862) );
  nand2_1 U15604 ( .A(n16223), .B(n16224), .Y(n16221) );
  o22ai_1 U15605 ( .A1(n16225), .A2(n16226), .B1(n16227), .B2(n16228), .Y(
        n16220) );
  nor2_1 U15606 ( .A(n16229), .B(n16224), .Y(n16227) );
  inv_1 U15607 ( .A(n16224), .Y(n16225) );
  o22ai_1 U15608 ( .A1(n771), .A2(n11211), .B1(n11213), .B2(n16230), .Y(n10305) );
  xor2_1 U15609 ( .A(n16231), .B(n16232), .X(n16230) );
  xor2_1 U15610 ( .A(n16233), .B(n16234), .X(n16232) );
  xor2_1 U15611 ( .A(n11249), .B(n11414), .X(n16231) );
  inv_1 U15612 ( .A(n23941), .Y(n11249) );
  mux2i_1 U15613 ( .A0(n16235), .A1(n16236), .S(n11213), .Y(n10304) );
  a22oi_1 U15614 ( .A1(n16206), .A2(n24054), .B1(n15718), .B2(n24048), .Y(
        n11213) );
  a211oi_1 U15615 ( .A1(n771), .A2(n16237), .B1(n11211), .C1(n11461), .Y(
        n16236) );
  xor2_1 U15616 ( .A(n16238), .B(n16239), .X(n16235) );
  xor2_1 U15617 ( .A(n23942), .B(n16240), .X(n16239) );
  inv_1 U15618 ( .A(n16241), .Y(n16238) );
  o32ai_1 U15619 ( .A1(n11480), .A2(n779), .A3(n11355), .B1(n16242), .B2(
        n11482), .Y(n10303) );
  xor2_1 U15620 ( .A(n16243), .B(n16244), .X(n16242) );
  xor2_1 U15621 ( .A(n16245), .B(n16246), .X(n16244) );
  xnor2_1 U15622 ( .A(n16247), .B(n16248), .Y(n16243) );
  o22ai_1 U15623 ( .A1(n16249), .A2(n16250), .B1(n16251), .B2(n16252), .Y(
        n10302) );
  xor2_1 U15624 ( .A(n16253), .B(n16254), .X(n16251) );
  xor2_1 U15625 ( .A(n20742), .B(n23740), .X(n16254) );
  or2_0 U15626 ( .A(n16255), .B(n20744), .X(n16253) );
  xor2_1 U15627 ( .A(n16256), .B(n16257), .X(n16250) );
  xor2_1 U15628 ( .A(n16258), .B(n16259), .X(n16257) );
  xor2_1 U15629 ( .A(n11489), .B(n40), .X(n16256) );
  o22ai_1 U15630 ( .A1(n16013), .A2(n16249), .B1(n16255), .B2(n16252), .Y(
        n10301) );
  o32ai_1 U15631 ( .A1(n16260), .A2(n12505), .A3(n16252), .B1(n16249), .B2(
        n16261), .Y(n10300) );
  xor2_1 U15632 ( .A(n16262), .B(n16263), .X(n16261) );
  nand2_1 U15633 ( .A(n16264), .B(n16265), .Y(n16263) );
  nand2_1 U15634 ( .A(n16266), .B(n16249), .Y(n16252) );
  xor2_1 U15635 ( .A(n20742), .B(n20744), .X(n16260) );
  nand2_1 U15636 ( .A(n16267), .B(n16268), .Y(n10299) );
  mux2i_1 U15637 ( .A0(n16269), .A1(n16270), .S(n16271), .Y(n16267) );
  xor2_1 U15638 ( .A(n16272), .B(n16273), .X(n16270) );
  xor2_1 U15639 ( .A(n16274), .B(n16275), .X(n16273) );
  xor2_1 U15640 ( .A(n16276), .B(n16277), .X(n16272) );
  xor2_1 U15641 ( .A(n16278), .B(n16279), .X(n16269) );
  nand2_1 U15642 ( .A(n23741), .B(n16280), .Y(n16279) );
  o22ai_1 U15643 ( .A1(n23760), .A2(n16281), .B1(n16282), .B2(n16283), .Y(
        n10298) );
  xor2_1 U15644 ( .A(n16284), .B(n16285), .X(n16283) );
  nor2_1 U15645 ( .A(n16286), .B(n16287), .Y(n16285) );
  xor2_1 U15646 ( .A(n16288), .B(n11159), .X(n16287) );
  nand2_1 U15647 ( .A(n16289), .B(n16268), .Y(n10297) );
  mux2i_1 U15648 ( .A0(n16290), .A1(n15953), .S(n16271), .Y(n16289) );
  nand2_1 U15649 ( .A(inData[22]), .B(n16291), .Y(n16290) );
  xor2_1 U15650 ( .A(n23741), .B(n23728), .X(n16291) );
  o32ai_1 U15651 ( .A1(n16292), .A2(n12826), .A3(n16281), .B1(n23951), .B2(
        n16282), .Y(n10296) );
  xor2_1 U15652 ( .A(n23741), .B(n2029), .X(n16292) );
  o32ai_1 U15653 ( .A1(n16281), .A2(n16293), .A3(n10679), .B1(n16282), .B2(
        n16294), .Y(n10295) );
  xor2_1 U15654 ( .A(n16295), .B(n16296), .X(n16294) );
  xnor2_1 U15655 ( .A(n23728), .B(n16297), .Y(n16296) );
  inv_1 U15656 ( .A(n12485), .Y(n16293) );
  mux2i_1 U15657 ( .A0(n15955), .A1(n16298), .S(n16282), .Y(n10294) );
  nor2_1 U15658 ( .A(n12570), .B(n16281), .Y(n16298) );
  nand2_1 U15659 ( .A(n16299), .B(n16300), .Y(n10293) );
  mux2i_1 U15660 ( .A0(n16301), .A1(n16302), .S(n16303), .Y(n16299) );
  xnor2_1 U15661 ( .A(n16304), .B(n16305), .Y(n16302) );
  xor2_1 U15662 ( .A(n16306), .B(n16307), .X(n16305) );
  nand2_1 U15663 ( .A(n16308), .B(inData[18]), .Y(n16301) );
  xor2_1 U15664 ( .A(n16309), .B(n16310), .X(n16308) );
  mux2i_1 U15665 ( .A0(n16311), .A1(n16312), .S(n16303), .Y(n10292) );
  xor2_1 U15666 ( .A(n16313), .B(n16314), .X(n16312) );
  xor2_1 U15667 ( .A(n16315), .B(n23737), .X(n16313) );
  nand3_1 U15668 ( .A(n16316), .B(n16317), .C(n16318), .Y(n16311) );
  a21oi_1 U15669 ( .A1(n16310), .A2(n40), .B1(n10675), .Y(n16318) );
  nor2_1 U15670 ( .A(n23738), .B(n23693), .Y(n16310) );
  o21ai_0 U15671 ( .A1(n23738), .A2(n16309), .B1(n23693), .Y(n16316) );
  inv_1 U15672 ( .A(n40), .Y(n16309) );
  nand2_1 U15673 ( .A(n16319), .B(n16300), .Y(n10291) );
  mux2i_1 U15674 ( .A0(n16320), .A1(n16321), .S(n16303), .Y(n16319) );
  xor2_1 U15675 ( .A(n16322), .B(n16323), .X(n16321) );
  xor2_1 U15676 ( .A(n16324), .B(n16325), .X(n16323) );
  xor2_1 U15677 ( .A(n10637), .B(n12959), .X(n16322) );
  nand2_1 U15678 ( .A(inData[26]), .B(n23763), .Y(n16320) );
  nand2_1 U15679 ( .A(n16326), .B(n16300), .Y(n10290) );
  mux2i_1 U15680 ( .A0(n23738), .A1(n23950), .S(n16303), .Y(n16326) );
  o32ai_1 U15681 ( .A1(n16327), .A2(n16328), .A3(n11775), .B1(n16329), .B2(
        n16330), .Y(n10289) );
  xor2_1 U15682 ( .A(n16331), .B(n16332), .X(n16330) );
  xor2_1 U15683 ( .A(n16333), .B(n12351), .X(n16328) );
  mux2i_1 U15684 ( .A0(n16334), .A1(n16335), .S(n16336), .Y(n10288) );
  nor3_1 U15685 ( .A(n11545), .B(n16337), .C(n16338), .Y(n16335) );
  xor2_1 U15686 ( .A(n23737), .B(n16339), .X(n16338) );
  xor2_1 U15687 ( .A(n16340), .B(n16341), .X(n16334) );
  xor2_1 U15688 ( .A(n23694), .B(n13031), .X(n16341) );
  xor2_1 U15689 ( .A(n16342), .B(n11554), .X(n16340) );
  mux2i_1 U15690 ( .A0(n12380), .A1(n16343), .S(n16336), .Y(n10287) );
  nor2_1 U15691 ( .A(n16337), .B(n16344), .Y(n16343) );
  xor2_1 U15692 ( .A(n20740), .B(n16345), .X(n16344) );
  inv_1 U15693 ( .A(n16346), .Y(n16337) );
  nand2_1 U15694 ( .A(n16347), .B(n16300), .Y(n10286) );
  mux2i_1 U15695 ( .A0(n23762), .A1(n16348), .S(n16303), .Y(n16347) );
  xor2_1 U15696 ( .A(n16349), .B(n16350), .X(n16348) );
  xor2_1 U15697 ( .A(n23720), .B(n16248), .X(n16349) );
  nand2_1 U15698 ( .A(n16351), .B(n16300), .Y(n10285) );
  or2_0 U15699 ( .A(n16317), .B(n16303), .X(n16300) );
  inv_1 U15700 ( .A(n16352), .Y(n16303) );
  nand2_1 U15701 ( .A(n16353), .B(n16354), .Y(n16317) );
  nand3_1 U15702 ( .A(n23893), .B(n14873), .C(n15978), .Y(n16354) );
  mux2_1 U15703 ( .A0(n23949), .A1(n16355), .S(n16352), .X(n16351) );
  nand4_1 U15704 ( .A(n16356), .B(n16005), .C(n16357), .D(n16358), .Y(n16352)
         );
  a21oi_1 U15705 ( .A1(n16359), .A2(n15457), .B1(n16360), .Y(n16358) );
  o21ai_0 U15706 ( .A1(n14873), .A2(n16361), .B1(n15887), .Y(n16359) );
  nand3_1 U15707 ( .A(n23893), .B(n23894), .C(n15978), .Y(n16357) );
  a211oi_1 U15708 ( .A1(n23762), .A2(n23737), .B1(n16345), .C1(n12699), .Y(
        n16355) );
  nor2_1 U15709 ( .A(n23762), .B(n23737), .Y(n16345) );
  o22ai_1 U15710 ( .A1(n16329), .A2(n16362), .B1(n16363), .B2(n16327), .Y(
        n10284) );
  xnor2_1 U15711 ( .A(n23694), .B(n16364), .Y(n16363) );
  nor2_1 U15712 ( .A(n12351), .B(n23736), .Y(n16364) );
  xor2_1 U15713 ( .A(n16365), .B(n16366), .X(n16362) );
  xor2_1 U15714 ( .A(n23750), .B(n12297), .X(n16366) );
  xor2_1 U15715 ( .A(n16367), .B(n10813), .X(n16365) );
  nand2_1 U15716 ( .A(n16368), .B(n16369), .Y(n10283) );
  mux2i_1 U15717 ( .A0(n16370), .A1(n16371), .S(n16329), .Y(n16368) );
  xor2_1 U15718 ( .A(n23765), .B(n12351), .X(n16371) );
  xor2_1 U15719 ( .A(n16372), .B(n16373), .X(n16370) );
  nor2_1 U15720 ( .A(n16374), .B(n16375), .Y(n16373) );
  inv_1 U15721 ( .A(n16376), .Y(n16374) );
  o32ai_1 U15722 ( .A1(n16377), .A2(n16378), .A3(n15993), .B1(n16379), .B2(
        n16336), .Y(n10282) );
  xor2_1 U15723 ( .A(n16380), .B(n16229), .X(n16379) );
  xor2_1 U15724 ( .A(n16381), .B(n23736), .X(n16380) );
  o22ai_1 U15725 ( .A1(n16382), .A2(n16336), .B1(n16383), .B2(n16377), .Y(
        n10281) );
  xor2_1 U15726 ( .A(n16378), .B(n23875), .X(n16383) );
  inv_1 U15727 ( .A(n23876), .Y(n16378) );
  xnor2_1 U15728 ( .A(n16384), .B(n16385), .Y(n16382) );
  nor2_1 U15729 ( .A(n16386), .B(n16387), .Y(n16385) );
  o22ai_1 U15730 ( .A1(n16336), .A2(n16388), .B1(n16389), .B2(n16377), .Y(
        n10280) );
  xor2_1 U15731 ( .A(n16390), .B(n43), .X(n16389) );
  nand2_1 U15732 ( .A(n23875), .B(n23876), .Y(n16390) );
  xor2_1 U15733 ( .A(n23876), .B(n16391), .X(n16388) );
  o32ai_1 U15734 ( .A1(n16377), .A2(n16392), .A3(n11775), .B1(n16393), .B2(
        n16336), .Y(n10279) );
  xor2_1 U15735 ( .A(n11779), .B(n16394), .X(n16393) );
  xor2_1 U15736 ( .A(n16395), .B(n16396), .X(n16394) );
  xor2_1 U15737 ( .A(n16397), .B(n23875), .X(n16392) );
  nand2_1 U15738 ( .A(n16346), .B(n16336), .Y(n16377) );
  nand4_1 U15739 ( .A(n15889), .B(n16398), .C(n16399), .D(n16400), .Y(n16336)
         );
  a221oi_1 U15740 ( .A1(n16401), .A2(n23894), .B1(n16402), .B2(n16403), .C1(
        n16404), .Y(n16400) );
  nor3_1 U15741 ( .A(n15457), .B(n16405), .C(n14873), .Y(n16404) );
  o21ai_0 U15742 ( .A1(n23895), .A2(n23892), .B1(n15888), .Y(n16403) );
  or2_0 U15743 ( .A(n15934), .B(n15951), .X(n15889) );
  o221ai_1 U15744 ( .A1(n23895), .A2(n16361), .B1(n23892), .B2(n16405), .C1(
        n15950), .Y(n16346) );
  inv_1 U15745 ( .A(n16406), .Y(n15950) );
  o211ai_1 U15746 ( .A1(n15934), .A2(n15887), .B1(n16005), .C1(n16398), .Y(
        n16406) );
  nand2_1 U15747 ( .A(n15963), .B(n16407), .Y(n16005) );
  o211ai_1 U15748 ( .A1(n16408), .A2(n16409), .B1(n23922), .C1(n16410), .Y(
        n10278) );
  mux2i_1 U15749 ( .A0(n16411), .A1(n16412), .S(n16413), .Y(n16410) );
  nor2_1 U15750 ( .A(n12584), .B(n16414), .Y(n16411) );
  xor2_1 U15751 ( .A(n16415), .B(n16413), .X(n16408) );
  o22ai_1 U15752 ( .A1(n12465), .A2(n10922), .B1(n16416), .B2(n10924), .Y(
        n10277) );
  xor2_1 U15753 ( .A(n16417), .B(n16418), .X(n16416) );
  xor2_1 U15754 ( .A(n16419), .B(n11131), .X(n16418) );
  xnor2_1 U15755 ( .A(n16420), .B(n16421), .Y(n16417) );
  nand2_1 U15756 ( .A(n16422), .B(n16423), .Y(n10276) );
  mux2i_1 U15757 ( .A0(n16424), .A1(n16425), .S(n16426), .Y(n16422) );
  or2_0 U15758 ( .A(n11355), .B(n12450), .X(n16425) );
  o22ai_1 U15759 ( .A1(n16427), .A2(n16428), .B1(n16429), .B2(n16430), .Y(
        n16424) );
  a21oi_1 U15760 ( .A1(n11130), .A2(n16431), .B1(n16427), .Y(n16430) );
  inv_1 U15761 ( .A(n28), .Y(n16431) );
  inv_1 U15762 ( .A(n16432), .Y(n16427) );
  nand2_1 U15763 ( .A(n16433), .B(n16423), .Y(n10275) );
  mux2i_1 U15764 ( .A0(n16434), .A1(n16435), .S(n16426), .Y(n16433) );
  nand2_1 U15765 ( .A(inData[24]), .B(n16436), .Y(n16435) );
  xor2_1 U15766 ( .A(n2047), .B(n16437), .X(n16436) );
  nor2_1 U15767 ( .A(n12450), .B(n23833), .Y(n16437) );
  o22ai_1 U15768 ( .A1(n16438), .A2(n16439), .B1(n16440), .B2(n16441), .Y(
        n16434) );
  and2_0 U15769 ( .A(n16442), .B(n16443), .X(n16440) );
  o32ai_1 U15770 ( .A1(n16444), .A2(n11330), .A3(n16445), .B1(n16426), .B2(
        n16446), .Y(n10274) );
  xor2_1 U15771 ( .A(n16447), .B(n16448), .X(n16446) );
  nand2_1 U15772 ( .A(n16449), .B(n16450), .Y(n16448) );
  xor2_1 U15773 ( .A(n23833), .B(n16451), .X(n16444) );
  nor2_1 U15774 ( .A(n12450), .B(n2047), .Y(n16451) );
  nand2_1 U15775 ( .A(n16452), .B(n16423), .Y(n10273) );
  mux2i_1 U15776 ( .A0(n16453), .A1(n16454), .S(n16426), .Y(n16452) );
  nand2_1 U15777 ( .A(inData[12]), .B(n28), .Y(n16454) );
  o22ai_1 U15778 ( .A1(n16455), .A2(n16445), .B1(n16426), .B2(n16456), .Y(
        n10272) );
  xor2_1 U15779 ( .A(n12725), .B(n16457), .X(n16456) );
  xor2_1 U15780 ( .A(n16458), .B(n23833), .X(n16457) );
  xor2_1 U15781 ( .A(n16459), .B(n12451), .X(n16455) );
  o22ai_1 U15782 ( .A1(n16460), .A2(n10922), .B1(n16461), .B2(n10924), .Y(
        n10271) );
  xor2_1 U15783 ( .A(n16462), .B(n16463), .X(n16461) );
  xor2_1 U15784 ( .A(n16464), .B(n16465), .X(n16463) );
  xor2_1 U15785 ( .A(n16466), .B(n16467), .X(n16462) );
  xor2_1 U15786 ( .A(n16468), .B(n16469), .X(n16460) );
  xor2_1 U15787 ( .A(outData[31]), .B(n23850), .X(n16469) );
  or2_0 U15788 ( .A(n12447), .B(n2046), .X(n16468) );
  o22ai_1 U15789 ( .A1(n23985), .A2(n16426), .B1(n16470), .B2(n16445), .Y(
        n10270) );
  xor2_1 U15790 ( .A(n16459), .B(n35), .X(n16470) );
  nand2_1 U15791 ( .A(n23843), .B(n12486), .Y(n16459) );
  nand2_1 U15792 ( .A(n16423), .B(n16445), .Y(n16426) );
  inv_1 U15793 ( .A(n16471), .Y(n16423) );
  o21ai_0 U15794 ( .A1(n23837), .A2(n16472), .B1(n16473), .Y(n16471) );
  nor2_1 U15795 ( .A(n10774), .B(n16474), .Y(n10269) );
  xor2_1 U15796 ( .A(n16475), .B(n16476), .X(n16474) );
  nor2_1 U15797 ( .A(n16477), .B(n16478), .Y(n16476) );
  inv_1 U15798 ( .A(n16479), .Y(n16477) );
  o32ai_1 U15799 ( .A1(n16480), .A2(n10923), .A3(n16473), .B1(n15445), .B2(
        n16481), .Y(n10268) );
  xor2_1 U15800 ( .A(n16482), .B(n16483), .X(n16481) );
  xor2_1 U15801 ( .A(n16484), .B(n27), .X(n16483) );
  inv_1 U15802 ( .A(n12583), .Y(n16480) );
  o32ai_1 U15803 ( .A1(n16485), .A2(n15993), .A3(n16473), .B1(n15990), .B2(
        n15445), .Y(n10267) );
  xnor2_1 U15804 ( .A(n37), .B(n16486), .Y(n16485) );
  nand2_1 U15805 ( .A(n26), .B(n16487), .Y(n16486) );
  mux2i_1 U15806 ( .A0(n16488), .A1(n16489), .S(n23836), .Y(n10266) );
  xor2_1 U15807 ( .A(n16490), .B(n16491), .X(n16489) );
  xor2_1 U15808 ( .A(n16492), .B(n16493), .X(n16491) );
  xor2_1 U15809 ( .A(n16494), .B(n16495), .X(n16490) );
  a211oi_1 U15810 ( .A1(n23754), .A2(n16492), .B1(n16473), .C1(n16496), .Y(
        n16488) );
  o32ai_1 U15811 ( .A1(n16497), .A2(n11134), .A3(n16473), .B1(n15445), .B2(
        n16498), .Y(n10265) );
  mux2i_1 U15812 ( .A0(n16499), .A1(n16500), .S(n12441), .Y(n16498) );
  xor2_1 U15813 ( .A(n16501), .B(n16502), .X(n16500) );
  xor2_1 U15814 ( .A(n16211), .B(n16502), .X(n16499) );
  xor2_1 U15815 ( .A(n16503), .B(n12939), .X(n16502) );
  xor2_1 U15816 ( .A(n27), .B(n16496), .X(n16497) );
  mux2i_1 U15817 ( .A0(n16504), .A1(n16505), .S(n23836), .Y(n10264) );
  xor2_1 U15818 ( .A(n16506), .B(n16507), .X(n16505) );
  xor2_1 U15819 ( .A(n12481), .B(n16508), .X(n16506) );
  nor3_1 U15820 ( .A(n16492), .B(n11330), .C(n16473), .Y(n16504) );
  o32ai_1 U15821 ( .A1(n16473), .A2(n16509), .A3(n11545), .B1(n16510), .B2(
        n15445), .Y(n10263) );
  xnor2_1 U15822 ( .A(n16496), .B(n12481), .Y(n16509) );
  nor2_1 U15823 ( .A(n16492), .B(n23754), .Y(n16496) );
  inv_1 U15824 ( .A(n23725), .Y(n16492) );
  nand2_1 U15825 ( .A(n15375), .B(n23837), .Y(n16473) );
  o22ai_1 U15826 ( .A1(n16511), .A2(n16512), .B1(n15445), .B2(n16513), .Y(
        n10262) );
  xor2_1 U15827 ( .A(n16514), .B(n16515), .X(n16513) );
  o21ai_0 U15828 ( .A1(n16516), .A2(n10640), .B1(n16517), .Y(n16515) );
  xor2_1 U15829 ( .A(n16518), .B(n16519), .X(n16511) );
  xor2_1 U15830 ( .A(n23753), .B(n2056), .X(n16519) );
  nand2_1 U15831 ( .A(n12480), .B(n23682), .Y(n16518) );
  o32ai_1 U15832 ( .A1(n16512), .A2(n16520), .A3(n11107), .B1(n16521), .B2(
        n15445), .Y(n10261) );
  xnor2_1 U15833 ( .A(n16522), .B(n16523), .Y(n16521) );
  xor2_1 U15834 ( .A(n16241), .B(n23730), .X(n16522) );
  o22ai_1 U15835 ( .A1(n16524), .A2(n15445), .B1(n2056), .B2(n16512), .Y(
        n10260) );
  nand2_1 U15836 ( .A(n16525), .B(n16526), .Y(n10259) );
  mux2i_1 U15837 ( .A0(n16527), .A1(n16528), .S(n16529), .Y(n16525) );
  nand2_1 U15838 ( .A(inData[2]), .B(n16530), .Y(n16528) );
  xor2_1 U15839 ( .A(n23757), .B(n23746), .X(n16530) );
  xor2_1 U15840 ( .A(n16531), .B(n16532), .X(n16527) );
  xor2_1 U15841 ( .A(n16533), .B(n16534), .X(n16532) );
  xor2_1 U15842 ( .A(n16535), .B(n12480), .X(n16531) );
  nand3_1 U15843 ( .A(n16536), .B(n16537), .C(n16538), .Y(n10258) );
  xnor2_1 U15844 ( .A(n2056), .B(n16539), .Y(n16538) );
  mux2i_1 U15845 ( .A0(n16540), .A1(n16541), .S(n23836), .Y(n16539) );
  xor2_1 U15846 ( .A(n16542), .B(n16543), .X(n16541) );
  o21ai_0 U15847 ( .A1(n10831), .A2(n10614), .B1(n15445), .Y(n16536) );
  nand2_1 U15848 ( .A(n16544), .B(n16526), .Y(n10257) );
  mux2i_1 U15849 ( .A0(n16545), .A1(n16546), .S(n16529), .Y(n16544) );
  xnor2_1 U15850 ( .A(n23745), .B(n16547), .Y(n16546) );
  nand2_1 U15851 ( .A(n23757), .B(n16548), .Y(n16547) );
  o32ai_1 U15852 ( .A1(n15898), .A2(n12475), .A3(n16537), .B1(n16529), .B2(
        n16549), .Y(n10256) );
  xor2_1 U15853 ( .A(n16550), .B(n16551), .X(n16549) );
  xor2_1 U15854 ( .A(n16552), .B(n23745), .X(n16551) );
  o22ai_1 U15855 ( .A1(n16529), .A2(n16553), .B1(n16537), .B2(n16554), .Y(
        n10255) );
  xor2_1 U15856 ( .A(n23757), .B(n23745), .X(n16554) );
  xor2_1 U15857 ( .A(n16555), .B(n16556), .X(n16553) );
  xor2_1 U15858 ( .A(n16216), .B(n16557), .X(n16556) );
  xor2_1 U15859 ( .A(n16548), .B(n11168), .X(n16555) );
  o22ai_1 U15860 ( .A1(n16558), .A2(n16537), .B1(n16559), .B2(n16529), .Y(
        n10254) );
  xor2_1 U15861 ( .A(n16560), .B(n16561), .X(n16559) );
  xor2_1 U15862 ( .A(n16562), .B(n23746), .X(n16560) );
  xor2_1 U15863 ( .A(n23733), .B(n16563), .X(n16558) );
  nand2_1 U15864 ( .A(n16564), .B(n16472), .Y(n10253) );
  mux2i_1 U15865 ( .A0(n16565), .A1(n16566), .S(n23836), .Y(n16564) );
  xor2_1 U15866 ( .A(n16567), .B(n16568), .X(n16566) );
  nand2_1 U15867 ( .A(inData[28]), .B(n23), .Y(n16565) );
  nand2_1 U15868 ( .A(n16569), .B(n16472), .Y(n10252) );
  mux2i_1 U15869 ( .A0(n16570), .A1(n12393), .S(n23836), .Y(n16569) );
  o211ai_1 U15870 ( .A1(n23), .A2(n16563), .B1(n16571), .C1(inData[30]), .Y(
        n16570) );
  nand2_1 U15871 ( .A(n16572), .B(n16472), .Y(n10251) );
  mux2i_1 U15872 ( .A0(n16573), .A1(n16574), .S(n23836), .Y(n16572) );
  xor2_1 U15873 ( .A(n11296), .B(n16575), .X(n16574) );
  xor2_1 U15874 ( .A(n22), .B(n16576), .X(n16575) );
  nand2_1 U15875 ( .A(n23683), .B(inData[20]), .Y(n16573) );
  nand3_1 U15876 ( .A(n16472), .B(n16577), .C(n16578), .Y(n10250) );
  mux2i_1 U15877 ( .A0(n11775), .A1(n10606), .S(n23836), .Y(n16578) );
  o22ai_1 U15878 ( .A1(n15445), .A2(n16579), .B1(n16580), .B2(n11545), .Y(
        n10249) );
  a22oi_1 U15879 ( .A1(n16581), .A2(n15375), .B1(n16582), .B2(n23756), .Y(
        n16580) );
  a21oi_1 U15880 ( .A1(n23756), .A2(n16577), .B1(n12441), .Y(n16581) );
  xor2_1 U15881 ( .A(n16583), .B(n16584), .X(n16579) );
  xor2_1 U15882 ( .A(n16585), .B(n23748), .X(n16584) );
  o21ai_0 U15883 ( .A1(n15445), .A2(n16586), .B1(n16587), .Y(n10248) );
  mux2i_1 U15884 ( .A0(n16582), .A1(n16588), .S(n23756), .Y(n16587) );
  a21oi_1 U15885 ( .A1(n12441), .A2(n16577), .B1(n16537), .Y(n16588) );
  nand2_1 U15886 ( .A(n23748), .B(n15445), .Y(n16577) );
  and3_1 U15887 ( .A(n15375), .B(n16589), .C(n12441), .X(n16582) );
  inv_1 U15888 ( .A(n16537), .Y(n15375) );
  xnor2_1 U15889 ( .A(n16590), .B(n16591), .Y(n16586) );
  nand2_1 U15890 ( .A(n16592), .B(n16593), .Y(n16590) );
  nand2_1 U15891 ( .A(n16594), .B(n16526), .Y(n10247) );
  nand2_1 U15892 ( .A(n16529), .B(n16537), .Y(n16526) );
  mux2i_1 U15893 ( .A0(n23958), .A1(n16595), .S(n16529), .Y(n16594) );
  nand2_1 U15894 ( .A(n23836), .B(n16445), .Y(n16529) );
  nand2_1 U15895 ( .A(n16596), .B(n23837), .Y(n16445) );
  xnor2_1 U15896 ( .A(n22), .B(n16571), .Y(n16595) );
  nand2_1 U15897 ( .A(n23), .B(n16563), .Y(n16571) );
  nand2_1 U15898 ( .A(n16597), .B(n16598), .Y(n10246) );
  mux2i_1 U15899 ( .A0(n16599), .A1(n16600), .S(n16601), .Y(n16597) );
  xor2_1 U15900 ( .A(n16602), .B(n16603), .X(n16600) );
  xor2_1 U15901 ( .A(n20741), .B(n23743), .X(n16603) );
  nor2_1 U15902 ( .A(n23742), .B(n16604), .Y(n16602) );
  inv_1 U15903 ( .A(n24), .Y(n16604) );
  xor2_1 U15904 ( .A(n16605), .B(n16606), .X(n16599) );
  xor2_1 U15905 ( .A(n10796), .B(n16607), .X(n16606) );
  mux2_1 U15906 ( .A0(n16608), .A1(n16609), .S(n12479), .X(n16605) );
  o32ai_1 U15907 ( .A1(n10831), .A2(n23742), .A3(n16610), .B1(n16611), .B2(
        n16601), .Y(n10245) );
  nand2_1 U15908 ( .A(n16612), .B(n16598), .Y(n10244) );
  mux2i_1 U15909 ( .A0(n16613), .A1(n16614), .S(n16601), .Y(n16612) );
  nand2_1 U15910 ( .A(inData[18]), .B(n16615), .Y(n16614) );
  xor2_1 U15911 ( .A(n20741), .B(n24), .X(n16615) );
  xnor2_1 U15912 ( .A(n16616), .B(n16617), .Y(n16613) );
  xor2_1 U15913 ( .A(n20741), .B(n11458), .X(n16616) );
  nand2_1 U15914 ( .A(n16618), .B(n16598), .Y(n10243) );
  nand2_1 U15915 ( .A(n16610), .B(n16601), .Y(n16598) );
  mux2i_1 U15916 ( .A0(n16619), .A1(n16620), .S(n16601), .Y(n16618) );
  xor2_1 U15917 ( .A(n16621), .B(n12516), .X(n16620) );
  xor2_1 U15918 ( .A(n16622), .B(n16623), .X(n16619) );
  xor2_1 U15919 ( .A(n16624), .B(n16625), .X(n16623) );
  xor2_1 U15920 ( .A(n16626), .B(n16627), .X(n16622) );
  o32ai_1 U15921 ( .A1(n16628), .A2(n11355), .A3(n16512), .B1(n15931), .B2(
        n15445), .Y(n10242) );
  o21ai_0 U15922 ( .A1(n20743), .A2(n16629), .B1(n16621), .Y(n16628) );
  o32ai_1 U15923 ( .A1(n11175), .A2(n16610), .A3(n16630), .B1(n23948), .B2(
        n16601), .Y(n10241) );
  xor2_1 U15924 ( .A(n16621), .B(n23730), .X(n16630) );
  nand2_1 U15925 ( .A(n20743), .B(n16629), .Y(n16621) );
  o32ai_1 U15926 ( .A1(n16512), .A2(n23758), .A3(n12699), .B1(n15445), .B2(
        n16631), .Y(n10240) );
  xnor2_1 U15927 ( .A(n16632), .B(n16633), .Y(n16631) );
  or2_0 U15928 ( .A(n16472), .B(n10614), .X(n16512) );
  nand2_1 U15929 ( .A(n15435), .B(n15445), .Y(n16472) );
  inv_1 U15930 ( .A(n23838), .Y(n15435) );
  o32ai_1 U15931 ( .A1(n10642), .A2(n16610), .A3(n10923), .B1(n16634), .B2(
        n16601), .Y(n10239) );
  xor2_1 U15932 ( .A(n16635), .B(n16636), .X(n16634) );
  xor2_1 U15933 ( .A(n10928), .B(n16637), .X(n16636) );
  xor2_1 U15934 ( .A(n16638), .B(n23742), .X(n16635) );
  nor2_1 U15935 ( .A(n16596), .B(n16639), .Y(n16610) );
  nor2_1 U15936 ( .A(n15445), .B(n23838), .Y(n16596) );
  nor2_1 U15937 ( .A(n16640), .B(n12628), .Y(n10238) );
  xor2_1 U15938 ( .A(n16641), .B(n16642), .X(n16640) );
  xor2_1 U15939 ( .A(n12583), .B(n12297), .X(n16642) );
  xor2_1 U15940 ( .A(n16643), .B(n16644), .X(n16641) );
  nor2_1 U15941 ( .A(n12628), .B(n16645), .Y(n10237) );
  xor2_1 U15942 ( .A(n12705), .B(n16646), .X(n16645) );
  xnor2_1 U15943 ( .A(n16647), .B(n16487), .Y(n16646) );
  inv_1 U15944 ( .A(n23830), .Y(n16487) );
  inv_1 U15945 ( .A(n12636), .Y(n12628) );
  a21oi_1 U15946 ( .A1(n16601), .A2(n23838), .B1(n16282), .Y(n12636) );
  nand2_1 U15947 ( .A(n16648), .B(n12652), .Y(n10236) );
  mux2i_1 U15948 ( .A0(n16649), .A1(n16650), .S(n12655), .Y(n16648) );
  nand2_1 U15949 ( .A(inData[10]), .B(n12666), .Y(n16650) );
  xor2_1 U15950 ( .A(n16651), .B(n16652), .X(n16649) );
  xnor2_1 U15951 ( .A(n16653), .B(n16654), .Y(n16652) );
  xor2_1 U15952 ( .A(n24045), .B(n16655), .X(n16651) );
  nor2_1 U15953 ( .A(n16656), .B(n10774), .Y(n10235) );
  xor2_1 U15954 ( .A(n11136), .B(n16657), .X(n16656) );
  xor2_1 U15955 ( .A(n16658), .B(n16659), .X(n16657) );
  nand2_1 U15956 ( .A(n16660), .B(n11032), .Y(n10234) );
  mux2i_1 U15957 ( .A0(n16661), .A1(n16662), .S(n11035), .Y(n16660) );
  xor2_1 U15958 ( .A(n18), .B(n16663), .X(n16662) );
  nor2_1 U15959 ( .A(n12430), .B(n23848), .Y(n16663) );
  xor2_1 U15960 ( .A(n16664), .B(n16665), .X(n16661) );
  xor2_1 U15961 ( .A(n16666), .B(n16667), .X(n16665) );
  xor2_1 U15962 ( .A(n16668), .B(n16669), .X(n16664) );
  nand2_1 U15963 ( .A(n16670), .B(n23922), .Y(n10233) );
  xor2_1 U15964 ( .A(n16671), .B(n16672), .X(n16670) );
  xor2_1 U15965 ( .A(n16673), .B(n12686), .X(n16672) );
  xor2_1 U15966 ( .A(n16674), .B(n16675), .X(n16671) );
  nand2_1 U15967 ( .A(n16676), .B(n11032), .Y(n10232) );
  nand2_1 U15968 ( .A(n16677), .B(n11035), .Y(n11032) );
  mux2i_1 U15969 ( .A0(n16678), .A1(n16679), .S(n11035), .Y(n16676) );
  o211ai_1 U15970 ( .A1(n24056), .A2(n16680), .B1(n16681), .C1(n16682), .Y(
        n11035) );
  nand2_1 U15971 ( .A(n16683), .B(inData[28]), .Y(n16679) );
  xor2_1 U15972 ( .A(n16684), .B(n23877), .X(n16683) );
  or2_0 U15973 ( .A(n16685), .B(n20), .X(n16684) );
  o22ai_1 U15974 ( .A1(n11057), .A2(n16686), .B1(n16687), .B2(n16688), .Y(
        n16678) );
  nor2_1 U15975 ( .A(n11057), .B(n16689), .Y(n16688) );
  xor2_1 U15976 ( .A(n12968), .B(n16690), .X(n16689) );
  nand2_1 U15977 ( .A(n11503), .B(n16691), .Y(n10231) );
  xor2_1 U15978 ( .A(n16692), .B(n16693), .X(n16691) );
  xor2_1 U15979 ( .A(n16694), .B(n16695), .X(n16693) );
  xor2_1 U15980 ( .A(n24045), .B(n2046), .X(n16692) );
  nand2_1 U15981 ( .A(n16696), .B(n11503), .Y(n10230) );
  xor2_1 U15982 ( .A(n16697), .B(n16698), .X(n16696) );
  xor2_1 U15983 ( .A(n16699), .B(n23850), .X(n16697) );
  mux2i_1 U15984 ( .A0(n16700), .A1(n16701), .S(n12663), .Y(n10229) );
  and3_1 U15985 ( .A(n10663), .B(n11045), .C(n23789), .X(n16701) );
  xor2_1 U15986 ( .A(n16702), .B(n16703), .X(n16700) );
  xor2_1 U15987 ( .A(n16704), .B(n16705), .X(n16703) );
  xor2_1 U15988 ( .A(n16706), .B(n16707), .X(n16702) );
  nor2_1 U15989 ( .A(n16708), .B(n10833), .Y(n10228) );
  xor2_1 U15990 ( .A(n16709), .B(n16710), .X(n16708) );
  xor2_1 U15991 ( .A(n16711), .B(n12517), .X(n16709) );
  o32ai_1 U15992 ( .A1(n11066), .A2(n16712), .A3(n12699), .B1(n11068), .B2(
        n16713), .Y(n10227) );
  xor2_1 U15993 ( .A(n16714), .B(n16715), .X(n16713) );
  xor2_1 U15994 ( .A(n16716), .B(n23878), .X(n16715) );
  xor2_1 U15995 ( .A(n11078), .B(n12518), .X(n16712) );
  o22ai_1 U15996 ( .A1(n11068), .A2(n16717), .B1(n11066), .B2(n16718), .Y(
        n10226) );
  xor2_1 U15997 ( .A(n11091), .B(n11078), .X(n16718) );
  nand2_1 U15998 ( .A(n41), .B(n20747), .Y(n11078) );
  xor2_1 U15999 ( .A(n16719), .B(n16720), .X(n16717) );
  xor2_1 U16000 ( .A(n16721), .B(n23848), .X(n16720) );
  inv_1 U16001 ( .A(n16722), .Y(n10225) );
  a211oi_1 U16002 ( .A1(n16723), .A2(n20), .B1(n16724), .C1(n10833), .Y(n16722) );
  o32ai_1 U16003 ( .A1(n16327), .A2(n23840), .A3(n10923), .B1(n16329), .B2(
        n16725), .Y(n10224) );
  inv_1 U16004 ( .A(n16726), .Y(n16725) );
  o22ai_1 U16005 ( .A1(n10797), .A2(n10798), .B1(n10826), .B2(n10800), .Y(
        n16726) );
  xor2_1 U16006 ( .A(n23750), .B(n10826), .X(n10798) );
  xnor2_1 U16007 ( .A(n16727), .B(n11284), .Y(n10797) );
  o22ai_1 U16008 ( .A1(n10813), .A2(n16367), .B1(n16728), .B2(n10800), .Y(
        n16727) );
  inv_1 U16009 ( .A(n23750), .Y(n10800) );
  and2_0 U16010 ( .A(n16367), .B(n10813), .X(n16728) );
  o22ai_1 U16011 ( .A1(n16229), .A2(n16381), .B1(n16729), .B2(n16333), .Y(
        n16367) );
  and2_0 U16012 ( .A(n16381), .B(n16229), .X(n16729) );
  o22ai_1 U16013 ( .A1(n16730), .A2(n16731), .B1(n16732), .B2(n16733), .Y(
        n16381) );
  inv_1 U16014 ( .A(n43), .Y(n16733) );
  and2_0 U16015 ( .A(n16731), .B(n16730), .X(n16732) );
  inv_1 U16016 ( .A(inData[16]), .Y(n10923) );
  o32ai_1 U16017 ( .A1(n16734), .A2(n10681), .A3(n16327), .B1(n16329), .B2(
        n16735), .Y(n10223) );
  a21oi_1 U16018 ( .A1(n16372), .A2(n16376), .B1(n16375), .Y(n16735) );
  xor2_1 U16019 ( .A(n16736), .B(n16737), .X(n16375) );
  nand2_1 U16020 ( .A(n16339), .B(n10826), .Y(n16736) );
  nand2_1 U16021 ( .A(n23720), .B(n12380), .Y(n16376) );
  a21oi_1 U16022 ( .A1(n16738), .A2(n16384), .B1(n16386), .Y(n16372) );
  nor2_1 U16023 ( .A(n16739), .B(n23720), .Y(n16386) );
  mux2_1 U16024 ( .A0(n16740), .A1(n16741), .S(n16742), .X(n16384) );
  or2_0 U16025 ( .A(n16332), .B(n16743), .X(n16741) );
  xor2_1 U16026 ( .A(n16744), .B(n16339), .X(n16332) );
  o22ai_1 U16027 ( .A1(n23720), .A2(n16743), .B1(n16745), .B2(n16744), .Y(
        n16740) );
  nor2_1 U16028 ( .A(n16339), .B(n16331), .Y(n16745) );
  inv_1 U16029 ( .A(n23720), .Y(n16339) );
  inv_1 U16030 ( .A(n16331), .Y(n16743) );
  o22ai_1 U16031 ( .A1(n16248), .A2(n16350), .B1(n23720), .B2(n16746), .Y(
        n16331) );
  and2_0 U16032 ( .A(n16248), .B(n16350), .X(n16746) );
  xnor2_1 U16033 ( .A(n16747), .B(n24045), .Y(n16350) );
  o22ai_1 U16034 ( .A1(n11666), .A2(n16324), .B1(n16748), .B2(n10637), .Y(
        n16747) );
  and2_0 U16035 ( .A(n16324), .B(n11666), .X(n16748) );
  o22ai_1 U16036 ( .A1(n16259), .A2(n16258), .B1(n40), .B2(n16749), .Y(n16324)
         );
  and2_0 U16037 ( .A(n16258), .B(n16259), .X(n16749) );
  xor2_1 U16038 ( .A(n12929), .B(n16750), .X(n16258) );
  a21oi_1 U16039 ( .A1(n16262), .A2(n16264), .B1(n16751), .Y(n16259) );
  inv_1 U16040 ( .A(n16265), .Y(n16751) );
  nand2_1 U16041 ( .A(n20742), .B(n16752), .Y(n16265) );
  xnor2_1 U16042 ( .A(n16753), .B(n16754), .Y(n16264) );
  nor2_1 U16043 ( .A(n20742), .B(n16752), .Y(n16754) );
  o21ai_0 U16044 ( .A1(n16288), .A2(n16284), .B1(n16755), .Y(n16262) );
  inv_1 U16045 ( .A(n16286), .Y(n16755) );
  xor2_1 U16046 ( .A(n16756), .B(n16757), .X(n16286) );
  nand2_1 U16047 ( .A(n16758), .B(n16278), .Y(n16756) );
  o22ai_1 U16048 ( .A1(n16295), .A2(n16297), .B1(n23728), .B2(n16759), .Y(
        n16284) );
  and2_0 U16049 ( .A(n16297), .B(n16295), .X(n16759) );
  o22ai_1 U16050 ( .A1(n16760), .A2(n16609), .B1(n12479), .B2(n16761), .Y(
        n16297) );
  nor2_1 U16051 ( .A(n16608), .B(n16607), .Y(n16761) );
  xor2_1 U16052 ( .A(n16762), .B(n16763), .X(n16609) );
  inv_1 U16053 ( .A(n16607), .Y(n16760) );
  o22ai_1 U16054 ( .A1(n16617), .A2(n11458), .B1(n16764), .B2(n10642), .Y(
        n16607) );
  and2_0 U16055 ( .A(n11458), .B(n16617), .X(n16764) );
  mux2i_1 U16056 ( .A0(n16765), .A1(n16766), .S(n11742), .Y(n16617) );
  o21ai_0 U16057 ( .A1(n16767), .A2(n16633), .B1(n16768), .Y(n16766) );
  nor2_1 U16058 ( .A(n16233), .B(n12516), .Y(n16767) );
  or2_0 U16059 ( .A(n16632), .B(n16633), .X(n16765) );
  xnor2_1 U16060 ( .A(n16769), .B(n13307), .Y(n16633) );
  o22ai_1 U16061 ( .A1(n16241), .A2(n16523), .B1(n16770), .B2(n16771), .Y(
        n16769) );
  inv_1 U16062 ( .A(n23730), .Y(n16771) );
  and2_0 U16063 ( .A(n16241), .B(n16523), .X(n16770) );
  xor2_1 U16064 ( .A(n16772), .B(n16773), .X(n16523) );
  o22ai_1 U16065 ( .A1(n16533), .A2(n16774), .B1(n16775), .B2(n16540), .Y(
        n16772) );
  inv_1 U16066 ( .A(n12480), .Y(n16540) );
  nor2_1 U16067 ( .A(n16534), .B(n16776), .Y(n16775) );
  inv_1 U16068 ( .A(n16774), .Y(n16534) );
  inv_1 U16069 ( .A(n16776), .Y(n16533) );
  o21ai_0 U16070 ( .A1(n12475), .A2(n16216), .B1(n16777), .Y(n16776) );
  xor2_1 U16071 ( .A(n16778), .B(n13351), .X(n16777) );
  nand2_1 U16072 ( .A(n16557), .B(n16779), .Y(n16778) );
  xor2_1 U16073 ( .A(n11751), .B(n16780), .X(n16779) );
  nor2_1 U16074 ( .A(n16781), .B(n16548), .Y(n16780) );
  inv_1 U16075 ( .A(n12475), .Y(n16548) );
  mux2_1 U16076 ( .A0(n16782), .A1(n16783), .S(n11520), .X(n16557) );
  nand2_1 U16077 ( .A(n16568), .B(n16784), .Y(n16783) );
  xor2_1 U16078 ( .A(n16785), .B(n23733), .X(n16568) );
  o22ai_1 U16079 ( .A1(n16567), .A2(n16785), .B1(n23733), .B2(n16786), .Y(
        n16782) );
  and2_0 U16080 ( .A(n16785), .B(n16567), .X(n16786) );
  inv_1 U16081 ( .A(n16784), .Y(n16567) );
  o22ai_1 U16082 ( .A1(n16576), .A2(n11296), .B1(n22), .B2(n16787), .Y(n16784)
         );
  nor2_1 U16083 ( .A(n16788), .B(n16789), .Y(n16787) );
  inv_1 U16084 ( .A(n16789), .Y(n16576) );
  o22ai_1 U16085 ( .A1(n16501), .A2(n16503), .B1(n12441), .B2(n16790), .Y(
        n16789) );
  and2_0 U16086 ( .A(n16503), .B(n16791), .X(n16790) );
  o22ai_1 U16087 ( .A1(n16495), .A2(n16792), .B1(n23725), .B2(n16793), .Y(
        n16503) );
  nor2_1 U16088 ( .A(n12519), .B(n16494), .Y(n16793) );
  inv_1 U16089 ( .A(n16494), .Y(n16792) );
  o22ai_1 U16090 ( .A1(n16644), .A2(n16643), .B1(n12583), .B2(n16794), .Y(
        n16494) );
  nor2_1 U16091 ( .A(n11155), .B(n16795), .Y(n16794) );
  inv_1 U16092 ( .A(n16795), .Y(n16644) );
  o21ai_0 U16093 ( .A1(n12635), .A2(n12632), .B1(n12633), .Y(n16795) );
  nand3_1 U16094 ( .A(n16450), .B(n16796), .C(n37), .Y(n12633) );
  a21oi_1 U16095 ( .A1(n16450), .A2(n16796), .B1(n37), .Y(n12635) );
  nand2_1 U16096 ( .A(n16449), .B(n16447), .Y(n16796) );
  nand2_1 U16097 ( .A(n16439), .B(n16442), .Y(n16447) );
  inv_1 U16098 ( .A(n16438), .Y(n16442) );
  nor2_1 U16099 ( .A(n11347), .B(n12450), .Y(n16438) );
  nand2_1 U16100 ( .A(n16443), .B(n16441), .Y(n16439) );
  o21ai_0 U16101 ( .A1(n16475), .A2(n16478), .B1(n16479), .Y(n16441) );
  nand2_1 U16102 ( .A(n12451), .B(n11548), .Y(n16479) );
  xor2_1 U16103 ( .A(n12968), .B(n16797), .X(n16478) );
  nor2_1 U16104 ( .A(n12451), .B(n11548), .Y(n16797) );
  a21oi_1 U16105 ( .A1(n12436), .A2(n12434), .B1(n12437), .Y(n16475) );
  xor2_1 U16106 ( .A(n11414), .B(n16798), .X(n12437) );
  nor2_1 U16107 ( .A(n16799), .B(n16800), .Y(n16798) );
  xnor2_1 U16108 ( .A(n16801), .B(n16802), .Y(n12434) );
  a21oi_1 U16109 ( .A1(n34), .A2(n16202), .B1(n16203), .Y(n16802) );
  nor2_1 U16110 ( .A(n16803), .B(n16804), .Y(n16203) );
  nand2_1 U16111 ( .A(n16804), .B(n16803), .Y(n16202) );
  o22ai_1 U16112 ( .A1(n16196), .A2(n16805), .B1(n12586), .B2(n16806), .Y(
        n16803) );
  nor2_1 U16113 ( .A(n16195), .B(n16197), .Y(n16806) );
  inv_1 U16114 ( .A(n16195), .Y(n16805) );
  a22oi_1 U16115 ( .A1(n10779), .A2(n10777), .B1(n16807), .B2(n23829), .Y(
        n16195) );
  or2_0 U16116 ( .A(n10777), .B(n10779), .X(n16807) );
  o22ai_1 U16117 ( .A1(n11779), .A2(n16396), .B1(n16808), .B2(n16395), .Y(
        n10779) );
  inv_1 U16118 ( .A(n36), .Y(n16395) );
  and2_0 U16119 ( .A(n16396), .B(n11779), .X(n16808) );
  nand3_1 U16120 ( .A(n16809), .B(n16810), .C(n16811), .Y(n16396) );
  xor2_1 U16121 ( .A(n12649), .B(n16812), .X(n16811) );
  nor3_1 U16122 ( .A(n16813), .B(n16814), .C(n16815), .Y(n16812) );
  mux2i_1 U16123 ( .A0(n16816), .A1(n16817), .S(n16818), .Y(n16815) );
  nor2_1 U16124 ( .A(n16819), .B(n16820), .Y(n16817) );
  mux2i_1 U16125 ( .A0(n16821), .A1(n16822), .S(n16823), .Y(n16820) );
  nand2_1 U16126 ( .A(n16822), .B(n16824), .Y(n16821) );
  a21oi_1 U16127 ( .A1(n16825), .A2(n16826), .B1(n24019), .Y(n16819) );
  mux2i_1 U16128 ( .A0(n16827), .A1(n16822), .S(n16823), .Y(n16816) );
  nor2_1 U16129 ( .A(n16828), .B(n16822), .Y(n16827) );
  xor2_1 U16130 ( .A(n16829), .B(n24019), .X(n16822) );
  xor2_1 U16131 ( .A(n16830), .B(n16831), .X(n16814) );
  xor2_1 U16132 ( .A(n16832), .B(n16833), .X(n16831) );
  nand2_1 U16133 ( .A(n16834), .B(n16835), .Y(n16830) );
  o32ai_1 U16134 ( .A1(n16836), .A2(n16825), .A3(n16837), .B1(n16824), .B2(
        n11336), .Y(n16813) );
  xnor2_1 U16135 ( .A(n16838), .B(n16839), .Y(n16810) );
  nand2_1 U16136 ( .A(n16840), .B(n16841), .Y(n16839) );
  xor2_1 U16137 ( .A(n16275), .B(n16842), .X(n16809) );
  xor2_1 U16138 ( .A(n16197), .B(n16843), .X(n16196) );
  nand2_1 U16139 ( .A(n16844), .B(n16800), .Y(n12436) );
  inv_1 U16140 ( .A(n35), .Y(n16800) );
  xor2_1 U16141 ( .A(n16845), .B(n16799), .X(n16844) );
  nand2_1 U16142 ( .A(n12450), .B(n16846), .Y(n16443) );
  xor2_1 U16143 ( .A(n12968), .B(n11347), .X(n16846) );
  xor2_1 U16144 ( .A(n16843), .B(n16847), .X(n16449) );
  nor2_1 U16145 ( .A(n23828), .B(n12744), .Y(n16847) );
  xnor2_1 U16146 ( .A(n16848), .B(n16849), .Y(n16450) );
  and2_0 U16147 ( .A(n12744), .B(n23828), .X(n16849) );
  xor2_1 U16148 ( .A(n16850), .B(n16211), .X(n16501) );
  o21ai_0 U16149 ( .A1(n12516), .A2(n16233), .B1(n16768), .Y(n16632) );
  xor2_1 U16150 ( .A(n16851), .B(n12959), .X(n16768) );
  nand2_1 U16151 ( .A(n12516), .B(n16233), .Y(n16851) );
  xnor2_1 U16152 ( .A(n12821), .B(n16852), .Y(n16288) );
  nor2_1 U16153 ( .A(n16758), .B(n16278), .Y(n16852) );
  inv_1 U16154 ( .A(n2029), .Y(n16278) );
  inv_1 U16155 ( .A(n16387), .Y(n16738) );
  xor2_1 U16156 ( .A(n16853), .B(n12942), .X(n16387) );
  nand2_1 U16157 ( .A(n23720), .B(n16739), .Y(n16853) );
  o21ai_0 U16158 ( .A1(n15977), .A2(n16360), .B1(n16329), .Y(n16327) );
  inv_1 U16159 ( .A(n15983), .Y(n16360) );
  xor2_1 U16160 ( .A(n31), .B(n23840), .X(n16734) );
  nand2_1 U16161 ( .A(n16854), .B(n16369), .Y(n10222) );
  nand3_1 U16162 ( .A(n15983), .B(n15966), .C(n16329), .Y(n16369) );
  a211oi_1 U16163 ( .A1(n23892), .A2(n15938), .B1(n16004), .C1(n16855), .Y(
        n15983) );
  nor2_1 U16164 ( .A(n15939), .B(n15951), .Y(n16004) );
  mux2i_1 U16165 ( .A0(n16856), .A1(n16857), .S(n16329), .Y(n16854) );
  and4_1 U16166 ( .A(n16858), .B(n15982), .C(n16859), .D(n16860), .X(n16329)
         );
  a211oi_1 U16167 ( .A1(n15977), .A2(n15457), .B1(n15959), .C1(n16861), .Y(
        n16860) );
  a21oi_1 U16168 ( .A1(n16399), .A2(n16353), .B1(n15939), .Y(n16861) );
  o32ai_1 U16169 ( .A1(n15457), .A2(n15951), .A3(n15311), .B1(n14873), .B2(
        n15939), .Y(n15959) );
  nand2_1 U16170 ( .A(n23892), .B(n15457), .Y(n15939) );
  inv_1 U16171 ( .A(n15966), .Y(n15977) );
  nand3_1 U16172 ( .A(n23893), .B(n23894), .C(n24037), .Y(n15966) );
  nand3_1 U16173 ( .A(n24037), .B(n23893), .C(n15963), .Y(n16859) );
  nand2_1 U16174 ( .A(n15978), .B(n15958), .Y(n15982) );
  nand3_1 U16175 ( .A(n15934), .B(n15304), .C(n15891), .Y(n16858) );
  inv_1 U16176 ( .A(n15967), .Y(n15891) );
  nand2_1 U16177 ( .A(n15311), .B(n14873), .Y(n15967) );
  nand2_1 U16178 ( .A(inData[16]), .B(n16333), .Y(n16857) );
  inv_1 U16179 ( .A(n23736), .Y(n16333) );
  xor2_1 U16180 ( .A(n11755), .B(n16862), .X(n16856) );
  xor2_1 U16181 ( .A(n16731), .B(n43), .X(n16862) );
  o22ai_1 U16182 ( .A1(n16342), .A2(n16863), .B1(n23694), .B2(n16864), .Y(
        n16731) );
  and2_0 U16183 ( .A(n16342), .B(n16863), .X(n16864) );
  o22ai_1 U16184 ( .A1(n16314), .A2(n16315), .B1(n23737), .B2(n16865), .Y(
        n16342) );
  and2_0 U16185 ( .A(n16315), .B(n16314), .X(n16865) );
  o22ai_1 U16186 ( .A1(n16304), .A2(n16307), .B1(n16866), .B2(n16306), .Y(
        n16315) );
  inv_1 U16187 ( .A(n23738), .Y(n16306) );
  and2_0 U16188 ( .A(n16307), .B(n16304), .X(n16866) );
  xor2_1 U16189 ( .A(n16867), .B(n16868), .X(n16304) );
  o22ai_1 U16190 ( .A1(n16869), .A2(n16870), .B1(n16871), .B2(n16255), .Y(
        n16867) );
  nor2_1 U16191 ( .A(n16872), .B(n16873), .Y(n16871) );
  inv_1 U16192 ( .A(n16873), .Y(n16869) );
  nand2_1 U16193 ( .A(n16874), .B(n16268), .Y(n10221) );
  or2_0 U16194 ( .A(n16266), .B(n16271), .X(n16268) );
  o211ai_1 U16195 ( .A1(n23894), .A2(n15981), .B1(n16356), .C1(n15975), .Y(
        n16266) );
  inv_1 U16196 ( .A(n16855), .Y(n15975) );
  o21ai_0 U16197 ( .A1(n15934), .A2(n16399), .B1(n15952), .Y(n16855) );
  nand4_1 U16198 ( .A(n15963), .B(n24037), .C(n23894), .D(n15311), .Y(n15952)
         );
  inv_1 U16199 ( .A(n15888), .Y(n15963) );
  inv_1 U16200 ( .A(n15938), .Y(n16399) );
  nand2_1 U16201 ( .A(n16407), .B(n15457), .Y(n16356) );
  mux2i_1 U16202 ( .A0(n16875), .A1(n16876), .S(n16271), .Y(n16874) );
  inv_1 U16203 ( .A(n16249), .Y(n16271) );
  o211ai_1 U16204 ( .A1(n16405), .A2(n15888), .B1(n16002), .C1(n15890), .Y(
        n16249) );
  and4_1 U16205 ( .A(n16361), .B(n16398), .C(n15941), .D(n16877), .X(n15890)
         );
  a222oi_1 U16206 ( .A1(n15943), .A2(n15457), .B1(n23892), .B2(n16407), .C1(
        n16401), .C2(n14873), .Y(n16877) );
  inv_1 U16207 ( .A(n15981), .Y(n16401) );
  nand2_1 U16208 ( .A(n15978), .B(n15311), .Y(n15981) );
  inv_1 U16209 ( .A(n15934), .Y(n15978) );
  nand2_1 U16210 ( .A(n23895), .B(n15184), .Y(n15934) );
  inv_1 U16211 ( .A(n16353), .Y(n16407) );
  nand2_1 U16212 ( .A(n15958), .B(n14873), .Y(n16353) );
  inv_1 U16213 ( .A(n15887), .Y(n15943) );
  nand2_1 U16214 ( .A(n16402), .B(n15311), .Y(n15887) );
  inv_1 U16215 ( .A(n15935), .Y(n16402) );
  nand2_1 U16216 ( .A(n24037), .B(n15304), .Y(n15935) );
  nand2_1 U16217 ( .A(n24037), .B(n15892), .Y(n15941) );
  inv_1 U16218 ( .A(n15936), .Y(n15892) );
  nand3_1 U16219 ( .A(n15184), .B(n15457), .C(n15958), .Y(n15936) );
  inv_1 U16220 ( .A(n16405), .Y(n15958) );
  inv_1 U16221 ( .A(n23895), .Y(n15457) );
  inv_1 U16222 ( .A(n15965), .Y(n16398) );
  nor4_1 U16223 ( .A(n15311), .B(n15951), .C(n23892), .D(n23895), .Y(n15965)
         );
  nand3_1 U16224 ( .A(n15184), .B(n15311), .C(n23894), .Y(n16361) );
  inv_1 U16225 ( .A(n23893), .Y(n15311) );
  inv_1 U16226 ( .A(n23892), .Y(n15184) );
  nand2_1 U16227 ( .A(n15938), .B(n23895), .Y(n16002) );
  nor2_1 U16228 ( .A(n15951), .B(n23893), .Y(n15938) );
  nand2_1 U16229 ( .A(n23894), .B(n14873), .Y(n15951) );
  inv_1 U16230 ( .A(n24037), .Y(n14873) );
  nand2_1 U16231 ( .A(n23895), .B(n23892), .Y(n15888) );
  nand2_1 U16232 ( .A(n23893), .B(n15304), .Y(n16405) );
  inv_1 U16233 ( .A(n23894), .Y(n15304) );
  xor2_1 U16234 ( .A(n16872), .B(n16878), .X(n16876) );
  xor2_1 U16235 ( .A(n16255), .B(n16873), .X(n16878) );
  o21ai_0 U16236 ( .A1(n16277), .A2(n16274), .B1(n16879), .Y(n16873) );
  xor2_1 U16237 ( .A(n16880), .B(n16881), .X(n16879) );
  a21oi_1 U16238 ( .A1(n16277), .A2(n16274), .B1(n16276), .Y(n16881) );
  o22ai_1 U16239 ( .A1(n16882), .A2(n16883), .B1(n23741), .B2(n16884), .Y(
        n16276) );
  and2_0 U16240 ( .A(n16883), .B(n16882), .X(n16884) );
  inv_1 U16241 ( .A(n23740), .Y(n16274) );
  inv_1 U16242 ( .A(n12513), .Y(n16255) );
  nand2_1 U16243 ( .A(n20742), .B(inData[20]), .Y(n16875) );
  o32ai_1 U16244 ( .A1(n16885), .A2(n15993), .A3(n16281), .B1(n16282), .B2(
        n16886), .Y(n10220) );
  xor2_1 U16245 ( .A(n16887), .B(n16888), .X(n16886) );
  xor2_1 U16246 ( .A(n12890), .B(n23727), .X(n16888) );
  xnor2_1 U16247 ( .A(n12479), .B(n16889), .Y(n16885) );
  nand2_1 U16248 ( .A(n23759), .B(n23727), .Y(n16889) );
  o32ai_1 U16249 ( .A1(n16281), .A2(n16890), .A3(n11775), .B1(n16282), .B2(
        n16891), .Y(n10219) );
  xor2_1 U16250 ( .A(n16892), .B(n16893), .X(n16891) );
  xor2_1 U16251 ( .A(n23741), .B(n12942), .X(n16893) );
  xor2_1 U16252 ( .A(n16883), .B(n16882), .X(n16892) );
  o22ai_1 U16253 ( .A1(n16887), .A2(n16894), .B1(n16895), .B2(n12570), .Y(
        n16883) );
  inv_1 U16254 ( .A(n23727), .Y(n12570) );
  nor2_1 U16255 ( .A(n12890), .B(n16896), .Y(n16895) );
  inv_1 U16256 ( .A(n16887), .Y(n16896) );
  xor2_1 U16257 ( .A(n16897), .B(n16898), .X(n16887) );
  o22ai_1 U16258 ( .A1(n16637), .A2(n16638), .B1(n23742), .B2(n16899), .Y(
        n16897) );
  and2_0 U16259 ( .A(n16638), .B(n16637), .X(n16899) );
  o22ai_1 U16260 ( .A1(n12907), .A2(n16624), .B1(n16900), .B2(n16626), .Y(
        n16638) );
  inv_1 U16261 ( .A(n23743), .Y(n16626) );
  and2_0 U16262 ( .A(n16624), .B(n12907), .X(n16900) );
  xnor2_1 U16263 ( .A(n16901), .B(n16902), .Y(n16624) );
  o21ai_0 U16264 ( .A1(n16516), .A2(n10640), .B1(n16903), .Y(n16901) );
  xor2_1 U16265 ( .A(n16904), .B(n16905), .X(n16903) );
  nand2_1 U16266 ( .A(n16514), .B(n16517), .Y(n16905) );
  nand2_1 U16267 ( .A(n16516), .B(n10640), .Y(n16517) );
  o22ai_1 U16268 ( .A1(n16543), .A2(n16906), .B1(n2056), .B2(n16907), .Y(
        n16514) );
  nor2_1 U16269 ( .A(n16542), .B(n16908), .Y(n16907) );
  inv_1 U16270 ( .A(n16908), .Y(n16543) );
  o22ai_1 U16271 ( .A1(n16550), .A2(n16552), .B1(n23745), .B2(n16909), .Y(
        n16908) );
  and2_0 U16272 ( .A(n16552), .B(n16550), .X(n16909) );
  o22ai_1 U16273 ( .A1(n16561), .A2(n16910), .B1(n23746), .B2(n16911), .Y(
        n16552) );
  nor2_1 U16274 ( .A(n16562), .B(n16912), .Y(n16911) );
  inv_1 U16275 ( .A(n16562), .Y(n16910) );
  xor2_1 U16276 ( .A(n16913), .B(n16914), .X(n16562) );
  nand2_1 U16277 ( .A(n16915), .B(n16593), .Y(n16913) );
  nand2_1 U16278 ( .A(n16916), .B(n16563), .Y(n16593) );
  inv_1 U16279 ( .A(n23747), .Y(n16563) );
  xor2_1 U16280 ( .A(n10868), .B(n16917), .X(n16915) );
  nor2_1 U16281 ( .A(n16918), .B(n16591), .Y(n16917) );
  xnor2_1 U16282 ( .A(n16919), .B(n10920), .Y(n16591) );
  o22ai_1 U16283 ( .A1(n16920), .A2(n16921), .B1(n16922), .B2(n16589), .Y(
        n16919) );
  inv_1 U16284 ( .A(n23748), .Y(n16589) );
  nor2_1 U16285 ( .A(n16583), .B(n16585), .Y(n16922) );
  inv_1 U16286 ( .A(n16585), .Y(n16920) );
  o22ai_1 U16287 ( .A1(n16507), .A2(n16508), .B1(n12481), .B2(n16923), .Y(
        n16585) );
  and2_0 U16288 ( .A(n16508), .B(n16507), .X(n16923) );
  o22ai_1 U16289 ( .A1(n16482), .A2(n16484), .B1(n27), .B2(n16924), .Y(n16508)
         );
  and2_0 U16290 ( .A(n16484), .B(n16482), .X(n16924) );
  o22ai_1 U16291 ( .A1(n16925), .A2(n16647), .B1(n23830), .B2(n16926), .Y(
        n16484) );
  and2_0 U16292 ( .A(n16647), .B(n16925), .X(n16926) );
  o22ai_1 U16293 ( .A1(n12638), .A2(n12640), .B1(n16927), .B2(n16928), .Y(
        n16647) );
  inv_1 U16294 ( .A(n23831), .Y(n16928) );
  nor2_1 U16295 ( .A(n12715), .B(n16929), .Y(n16927) );
  inv_1 U16296 ( .A(n12638), .Y(n16929) );
  xor2_1 U16297 ( .A(n16930), .B(n16931), .X(n12638) );
  nand2_1 U16298 ( .A(n16932), .B(n16432), .Y(n16930) );
  nand2_1 U16299 ( .A(n28), .B(n16933), .Y(n16432) );
  xor2_1 U16300 ( .A(n16934), .B(n16428), .X(n16932) );
  o21ai_0 U16301 ( .A1(n28), .A2(n16933), .B1(n16429), .Y(n16428) );
  inv_1 U16302 ( .A(n16935), .Y(n16429) );
  o22ai_1 U16303 ( .A1(n12725), .A2(n16458), .B1(n16936), .B2(n10645), .Y(
        n16935) );
  and2_0 U16304 ( .A(n16458), .B(n12725), .X(n16936) );
  o22ai_1 U16305 ( .A1(n16937), .A2(n16938), .B1(n16939), .B2(n16658), .Y(
        n16458) );
  inv_1 U16306 ( .A(n12486), .Y(n16658) );
  nor2_1 U16307 ( .A(n11136), .B(n16659), .Y(n16939) );
  inv_1 U16308 ( .A(n16659), .Y(n16937) );
  o22ai_1 U16309 ( .A1(n16940), .A2(n12444), .B1(n1144), .B2(n16941), .Y(
        n16659) );
  and2_0 U16310 ( .A(n12444), .B(n16940), .X(n16941) );
  o22ai_1 U16311 ( .A1(n12731), .A2(n16942), .B1(n16943), .B2(n16673), .Y(
        n12444) );
  inv_1 U16312 ( .A(n39), .Y(n16673) );
  nor2_1 U16313 ( .A(n16675), .B(n16674), .Y(n16943) );
  inv_1 U16314 ( .A(n16942), .Y(n16675) );
  o21ai_0 U16315 ( .A1(n16414), .A2(n16409), .B1(n16944), .Y(n16942) );
  xor2_1 U16316 ( .A(n12726), .B(n16945), .X(n16944) );
  or2_0 U16317 ( .A(n16413), .B(n16412), .X(n16945) );
  nor2_1 U16318 ( .A(n16415), .B(n12584), .Y(n16412) );
  inv_1 U16319 ( .A(n16946), .Y(n16413) );
  o21ai_0 U16320 ( .A1(n10789), .A2(n10786), .B1(n10788), .Y(n16946) );
  nand2_1 U16321 ( .A(n23686), .B(n11120), .Y(n10788) );
  nand2_1 U16322 ( .A(n23876), .B(n16947), .Y(n10786) );
  nor2_1 U16323 ( .A(n11120), .B(n23686), .Y(n10789) );
  inv_1 U16324 ( .A(n12584), .Y(n16409) );
  inv_1 U16325 ( .A(n16592), .Y(n16918) );
  nand2_1 U16326 ( .A(n23747), .B(n16948), .Y(n16592) );
  and2_0 U16327 ( .A(n10614), .B(n16601), .X(n16282) );
  nand2_1 U16328 ( .A(n23838), .B(n23836), .Y(n16601) );
  inv_1 U16329 ( .A(inData[2]), .Y(n11775) );
  xor2_1 U16330 ( .A(n16949), .B(n23759), .X(n16890) );
  nand2_1 U16331 ( .A(n12479), .B(n23727), .Y(n16949) );
  inv_1 U16332 ( .A(n16639), .Y(n16281) );
  nor2_1 U16333 ( .A(n16537), .B(n23837), .Y(n16639) );
  nand2_1 U16334 ( .A(n23838), .B(n15445), .Y(n16537) );
  inv_1 U16335 ( .A(n23836), .Y(n15445) );
  nand2_1 U16336 ( .A(n16950), .B(n16951), .Y(n10218) );
  mux2i_1 U16337 ( .A0(n16952), .A1(n16953), .S(n11402), .Y(n16950) );
  nand2_1 U16338 ( .A(n16954), .B(inData[0]), .Y(n16953) );
  xnor2_1 U16339 ( .A(n11461), .B(n12484), .Y(n16954) );
  nor2_1 U16340 ( .A(n16237), .B(n771), .Y(n11461) );
  inv_1 U16341 ( .A(n67), .Y(n16237) );
  xor2_1 U16342 ( .A(n16955), .B(n16956), .X(n16952) );
  xor2_1 U16343 ( .A(n16762), .B(n769), .X(n16956) );
  nand2_1 U16344 ( .A(n16957), .B(n16951), .Y(n10217) );
  mux2i_1 U16345 ( .A0(n16958), .A1(n16959), .S(n11402), .Y(n16957) );
  xor2_1 U16346 ( .A(n16752), .B(n16960), .X(n16958) );
  xor2_1 U16347 ( .A(n16961), .B(n69), .X(n16960) );
  nand2_1 U16348 ( .A(n16962), .B(n16951), .Y(n10216) );
  mux2i_1 U16349 ( .A0(n16963), .A1(n16964), .S(n11402), .Y(n16962) );
  nand2_1 U16350 ( .A(n16965), .B(inData[8]), .Y(n16964) );
  xor2_1 U16351 ( .A(n16966), .B(n68), .X(n16965) );
  xor2_1 U16352 ( .A(n16967), .B(n16968), .X(n16963) );
  xor2_1 U16353 ( .A(n16969), .B(n16295), .X(n16968) );
  xor2_1 U16354 ( .A(n11394), .B(n16801), .X(n16967) );
  nand2_1 U16355 ( .A(n16970), .B(n16971), .Y(n10215) );
  mux2i_1 U16356 ( .A0(n16972), .A1(n16973), .S(n16974), .Y(n16970) );
  nand2_1 U16357 ( .A(inData[4]), .B(n23697), .Y(n16973) );
  xor2_1 U16358 ( .A(n16975), .B(n16976), .X(n16972) );
  xor2_1 U16359 ( .A(n10634), .B(n16977), .X(n16976) );
  o32ai_1 U16360 ( .A1(n16978), .A2(n16979), .A3(n11330), .B1(n16974), .B2(
        n16980), .Y(n10214) );
  xor2_1 U16361 ( .A(n16981), .B(n16982), .X(n16980) );
  inv_1 U16362 ( .A(inData[4]), .Y(n11330) );
  xor2_1 U16363 ( .A(n16983), .B(n16984), .X(n16978) );
  nand2_1 U16364 ( .A(n23697), .B(n16985), .Y(n16984) );
  o32ai_1 U16365 ( .A1(n12866), .A2(n10), .A3(n12826), .B1(n12863), .B2(n16986), .Y(n10213) );
  xor2_1 U16366 ( .A(n16987), .B(n16988), .X(n16986) );
  xor2_1 U16367 ( .A(n16989), .B(n16990), .X(n16988) );
  o22ai_1 U16368 ( .A1(n23884), .A2(n16991), .B1(n16992), .B2(n12887), .Y(
        n10212) );
  xor2_1 U16369 ( .A(n16993), .B(n16994), .X(n16992) );
  xor2_1 U16370 ( .A(n12372), .B(n16995), .X(n16994) );
  xor2_1 U16371 ( .A(n16872), .B(n16996), .X(n16993) );
  o22ai_1 U16372 ( .A1(n12887), .A2(n16997), .B1(n16998), .B2(n16991), .Y(
        n10211) );
  xor2_1 U16373 ( .A(n16999), .B(n12446), .X(n16998) );
  nand2_1 U16374 ( .A(n12445), .B(n17000), .Y(n16999) );
  xor2_1 U16375 ( .A(n17001), .B(n17002), .X(n16997) );
  a21oi_1 U16376 ( .A1(n17003), .A2(n17004), .B1(n17005), .Y(n17002) );
  o22ai_1 U16377 ( .A1(n12887), .A2(n17006), .B1(n17007), .B2(n16991), .Y(
        n10210) );
  nand2_1 U16378 ( .A(n12884), .B(n12887), .Y(n16991) );
  nand4_1 U16379 ( .A(n17008), .B(n17009), .C(n17010), .D(n15860), .Y(n12884)
         );
  o21ai_0 U16380 ( .A1(n15867), .A2(n17011), .B1(n24059), .Y(n17010) );
  nand2_1 U16381 ( .A(n11438), .B(n15867), .Y(n17009) );
  xnor2_1 U16382 ( .A(n12445), .B(n17012), .Y(n17007) );
  nor2_1 U16383 ( .A(n12446), .B(n23884), .Y(n17012) );
  xor2_1 U16384 ( .A(n17013), .B(n17014), .X(n17006) );
  o21ai_0 U16385 ( .A1(n17015), .A2(n12915), .B1(n17016), .Y(n12887) );
  a21oi_1 U16386 ( .A1(n15835), .A2(n24053), .B1(n11453), .Y(n17015) );
  o32ai_1 U16387 ( .A1(n12826), .A2(n17017), .A3(n11472), .B1(n11470), .B2(
        n17018), .Y(n10209) );
  xor2_1 U16388 ( .A(n17019), .B(n17020), .X(n17018) );
  a21oi_1 U16389 ( .A1(n17021), .A2(n16799), .B1(n17022), .Y(n17019) );
  o22ai_1 U16390 ( .A1(n11470), .A2(n17023), .B1(n11472), .B2(n17024), .Y(
        n10208) );
  o21ai_0 U16391 ( .A1(n12547), .A2(n12549), .B1(n11343), .Y(n17024) );
  nand2_1 U16392 ( .A(n12549), .B(n12547), .Y(n11343) );
  or2_0 U16393 ( .A(n16206), .B(n24054), .X(n11472) );
  xor2_1 U16394 ( .A(n17025), .B(n17026), .X(n17023) );
  xnor2_1 U16395 ( .A(n17027), .B(n16804), .Y(n17026) );
  xor2_1 U16396 ( .A(n16246), .B(n23925), .X(n17025) );
  nor2_1 U16397 ( .A(n15718), .B(n15870), .Y(n11470) );
  nand2_1 U16398 ( .A(n17028), .B(n23922), .Y(n10207) );
  xnor2_1 U16399 ( .A(n17029), .B(n17030), .Y(n17028) );
  xor2_1 U16400 ( .A(n17031), .B(n17032), .X(n17030) );
  or2_0 U16401 ( .A(n48), .B(n11558), .X(n10206) );
  nand2_1 U16402 ( .A(n23922), .B(n17033), .Y(n10205) );
  xor2_1 U16403 ( .A(n17034), .B(n17035), .X(n17033) );
  xor2_1 U16404 ( .A(n17036), .B(n17037), .X(n17035) );
  nand2_1 U16405 ( .A(n17038), .B(n23922), .Y(n10204) );
  xnor2_1 U16406 ( .A(n17039), .B(n17040), .Y(n17038) );
  xor2_1 U16407 ( .A(n17041), .B(n17042), .X(n17039) );
  nor2_1 U16408 ( .A(n17043), .B(n10774), .Y(n10203) );
  xnor2_1 U16409 ( .A(n17044), .B(n17045), .Y(n17043) );
  xor2_1 U16410 ( .A(n17046), .B(n17047), .X(n17045) );
  o32ai_1 U16411 ( .A1(n17048), .A2(n11415), .A3(n17049), .B1(n10924), .B2(
        n17050), .Y(n10202) );
  inv_1 U16412 ( .A(n65), .Y(n17050) );
  nand2_1 U16413 ( .A(n15795), .B(n11703), .Y(n10924) );
  a21oi_1 U16414 ( .A1(outData[21]), .A2(outData[19]), .B1(outData[20]), .Y(
        n17049) );
  nor2_1 U16415 ( .A(n12552), .B(n11495), .Y(n11415) );
  inv_1 U16416 ( .A(n11703), .Y(n11495) );
  inv_1 U16417 ( .A(n10922), .Y(n12552) );
  nand2_1 U16418 ( .A(n24062), .B(n12551), .Y(n10922) );
  o21ai_0 U16419 ( .A1(n17051), .A2(n12977), .B1(inData[2]), .Y(n17048) );
  o32ai_1 U16420 ( .A1(n17052), .A2(n17053), .A3(n17054), .B1(n17055), .B2(
        n17056), .Y(n10201) );
  xor2_1 U16421 ( .A(n17057), .B(n17058), .X(n17056) );
  a21oi_1 U16422 ( .A1(n17059), .A2(n17060), .B1(n17061), .Y(n17058) );
  o21ai_0 U16423 ( .A1(n23775), .A2(n20746), .B1(inData[28]), .Y(n17052) );
  o32ai_1 U16424 ( .A1(n10676), .A2(n17062), .A3(n11066), .B1(n17063), .B2(
        n11068), .Y(n10200) );
  xor2_1 U16425 ( .A(n17064), .B(n17065), .X(n17063) );
  xor2_1 U16426 ( .A(n17066), .B(n17067), .X(n17065) );
  xor2_1 U16427 ( .A(n17068), .B(n17069), .X(n17064) );
  xor2_1 U16428 ( .A(n17054), .B(n17070), .X(n17062) );
  o22ai_1 U16429 ( .A1(n17071), .A2(n11068), .B1(n17072), .B2(n11066), .Y(
        n10199) );
  o21ai_0 U16430 ( .A1(n17073), .A2(n17074), .B1(n11068), .Y(n11066) );
  inv_1 U16431 ( .A(n11075), .Y(n17073) );
  xor2_1 U16432 ( .A(n17054), .B(n17075), .X(n17072) );
  nor2_1 U16433 ( .A(n17076), .B(n10632), .Y(n17054) );
  nand2_1 U16434 ( .A(n16682), .B(n11075), .Y(n11068) );
  o21ai_0 U16435 ( .A1(n15714), .A2(n15789), .B1(n10613), .Y(n11075) );
  inv_1 U16436 ( .A(n15801), .Y(n15789) );
  inv_1 U16437 ( .A(n17077), .Y(n15714) );
  and3_1 U16438 ( .A(n11084), .B(n15740), .C(n17078), .X(n16682) );
  xnor2_1 U16439 ( .A(n17079), .B(n17080), .Y(n17071) );
  nand2_1 U16440 ( .A(n17081), .B(n17082), .Y(n17079) );
  o32ai_1 U16441 ( .A1(n17076), .A2(n17053), .A3(n11107), .B1(n17055), .B2(
        n17083), .Y(n10198) );
  xor2_1 U16442 ( .A(n17084), .B(n17085), .X(n17083) );
  xnor2_1 U16443 ( .A(n17086), .B(n17087), .Y(n17085) );
  xor2_1 U16444 ( .A(n11520), .B(n17088), .X(n17084) );
  mux2i_1 U16445 ( .A0(n17089), .A1(n17090), .S(n17055), .Y(n10197) );
  nor3_1 U16446 ( .A(n17091), .B(n17053), .C(n11107), .Y(n17090) );
  xor2_1 U16447 ( .A(n23779), .B(n23778), .X(n17091) );
  xor2_1 U16448 ( .A(n17092), .B(n17093), .X(n17089) );
  mux2i_1 U16449 ( .A0(n17094), .A1(n17095), .S(n17055), .Y(n10196) );
  nor3_1 U16450 ( .A(n17096), .B(n17053), .C(n15898), .Y(n17095) );
  xor2_1 U16451 ( .A(n23783), .B(n23779), .X(n17096) );
  xor2_1 U16452 ( .A(n17097), .B(n17098), .X(n17094) );
  nand2_1 U16453 ( .A(n17099), .B(n17100), .Y(n17098) );
  inv_1 U16454 ( .A(n17101), .Y(n17099) );
  o32ai_1 U16455 ( .A1(n17102), .A2(n17053), .A3(n12826), .B1(n17055), .B2(
        n17103), .Y(n10195) );
  xor2_1 U16456 ( .A(n17104), .B(n17105), .X(n17103) );
  xor2_1 U16457 ( .A(n17106), .B(n17107), .X(n17105) );
  xor2_1 U16458 ( .A(n10946), .B(n17108), .X(n17104) );
  inv_1 U16459 ( .A(inData[0]), .Y(n12826) );
  xnor2_1 U16460 ( .A(n23778), .B(n17109), .Y(n17102) );
  nand2_1 U16461 ( .A(n23784), .B(n23779), .Y(n17109) );
  o22ai_1 U16462 ( .A1(n17053), .A2(n10643), .B1(n17055), .B2(n17110), .Y(
        n10194) );
  xor2_1 U16463 ( .A(n17111), .B(n17112), .X(n17110) );
  o21ai_0 U16464 ( .A1(n17113), .A2(n17114), .B1(n17115), .Y(n17111) );
  nand3_1 U16465 ( .A(n17078), .B(n17116), .C(n17053), .Y(n17055) );
  inv_1 U16466 ( .A(n17117), .Y(n17078) );
  o21ai_0 U16467 ( .A1(n10613), .A2(n15827), .B1(n17118), .Y(n17117) );
  and3_1 U16468 ( .A(n16681), .B(n15865), .C(n17119), .X(n17053) );
  nand2_1 U16469 ( .A(n17120), .B(n11593), .Y(n10193) );
  mux2i_1 U16470 ( .A0(n17121), .A1(n17122), .S(n10819), .Y(n17120) );
  nand2_1 U16471 ( .A(inData[26]), .B(n11598), .Y(n17122) );
  inv_1 U16472 ( .A(n23799), .Y(n11598) );
  xor2_1 U16473 ( .A(n11727), .B(n17123), .X(n17121) );
  xor2_1 U16474 ( .A(n17124), .B(n16), .X(n17123) );
  mux2i_1 U16475 ( .A0(n17125), .A1(n17126), .S(n11087), .Y(n10192) );
  nor3_1 U16476 ( .A(n17127), .B(n16677), .C(n17128), .Y(n17126) );
  o21ai_0 U16477 ( .A1(n23796), .A2(n23766), .B1(inData[10]), .Y(n17127) );
  xor2_1 U16478 ( .A(n17129), .B(n17130), .X(n17125) );
  xor2_1 U16479 ( .A(n17131), .B(n17132), .X(n17130) );
  xor2_1 U16480 ( .A(n17070), .B(n17133), .X(n17129) );
  mux2i_1 U16481 ( .A0(n17134), .A1(n17135), .S(n11087), .Y(n10191) );
  nor3_1 U16482 ( .A(n17136), .B(n16677), .C(n11545), .Y(n17135) );
  xor2_1 U16483 ( .A(n23795), .B(n17128), .X(n17136) );
  xor2_1 U16484 ( .A(n17137), .B(n17138), .X(n17134) );
  xor2_1 U16485 ( .A(n17139), .B(n23774), .X(n17137) );
  o22ai_1 U16486 ( .A1(n11087), .A2(n17140), .B1(n11084), .B2(n17141), .Y(
        n10190) );
  xor2_1 U16487 ( .A(n23787), .B(n17128), .X(n17141) );
  nor2_1 U16488 ( .A(n17142), .B(n10625), .Y(n17128) );
  xor2_1 U16489 ( .A(n17143), .B(n17144), .X(n17140) );
  xor2_1 U16490 ( .A(n17145), .B(n17146), .X(n17144) );
  xor2_1 U16491 ( .A(n17076), .B(n12817), .X(n17143) );
  inv_1 U16492 ( .A(n23775), .Y(n17076) );
  o32ai_1 U16493 ( .A1(n15993), .A2(n10625), .A3(n11084), .B1(n11087), .B2(
        n17147), .Y(n10189) );
  xor2_1 U16494 ( .A(n17148), .B(n17149), .X(n17147) );
  o21ai_0 U16495 ( .A1(n17150), .A2(n10632), .B1(n17151), .Y(n17149) );
  xor2_1 U16496 ( .A(n17152), .B(n17153), .X(n17151) );
  inv_1 U16497 ( .A(inData[12]), .Y(n15993) );
  nand2_1 U16498 ( .A(n17154), .B(n12652), .Y(n10188) );
  mux2i_1 U16499 ( .A0(n17155), .A1(n17156), .S(n12655), .Y(n17154) );
  xor2_1 U16500 ( .A(n17157), .B(n17158), .X(n17156) );
  xor2_1 U16501 ( .A(n17159), .B(n17160), .X(n17155) );
  xor2_1 U16502 ( .A(n17161), .B(n17162), .X(n17159) );
  nand2_1 U16503 ( .A(n17163), .B(n12652), .Y(n10187) );
  nand2_1 U16504 ( .A(n11074), .B(n12655), .Y(n12652) );
  mux2i_1 U16505 ( .A0(n17164), .A1(n23781), .S(n12655), .Y(n17163) );
  xor2_1 U16506 ( .A(n17165), .B(n17166), .X(n17164) );
  xnor2_1 U16507 ( .A(n17167), .B(n17168), .Y(n17165) );
  mux2i_1 U16508 ( .A0(n17169), .A1(n17170), .S(n12655), .Y(n10186) );
  nand2_1 U16509 ( .A(n17171), .B(n17074), .Y(n17170) );
  xor2_1 U16510 ( .A(n23781), .B(n23696), .X(n17171) );
  xnor2_1 U16511 ( .A(n17172), .B(n17173), .Y(n17169) );
  xor2_1 U16512 ( .A(n17174), .B(n17175), .X(n17173) );
  nand2_1 U16513 ( .A(n17176), .B(n17177), .Y(n17175) );
  inv_1 U16514 ( .A(n17178), .Y(n17176) );
  mux2i_1 U16515 ( .A0(n17179), .A1(n17180), .S(n12655), .Y(n10185) );
  nand3_1 U16516 ( .A(n17119), .B(n15827), .C(n16677), .Y(n12655) );
  nand2_1 U16517 ( .A(n17181), .B(n17074), .Y(n17180) );
  xor2_1 U16518 ( .A(n23691), .B(n17158), .X(n17181) );
  nor2_1 U16519 ( .A(n23781), .B(n23696), .Y(n17158) );
  xor2_1 U16520 ( .A(n17182), .B(n17183), .X(n17179) );
  nand2_1 U16521 ( .A(n17184), .B(n16971), .Y(n10184) );
  mux2i_1 U16522 ( .A0(n17185), .A1(n17186), .S(n16974), .Y(n17184) );
  xor2_1 U16523 ( .A(n16985), .B(n23794), .X(n17186) );
  xor2_1 U16524 ( .A(n17187), .B(n17188), .X(n17185) );
  xor2_1 U16525 ( .A(n16848), .B(n17189), .X(n17188) );
  nand2_1 U16526 ( .A(n17190), .B(n16971), .Y(n10183) );
  nand2_1 U16527 ( .A(n16974), .B(n16979), .Y(n16971) );
  mux2i_1 U16528 ( .A0(n17191), .A1(n17192), .S(n16974), .Y(n17190) );
  xor2_1 U16529 ( .A(n12544), .B(n16985), .X(n17192) );
  xnor2_1 U16530 ( .A(n17193), .B(n17194), .Y(n17191) );
  xor2_1 U16531 ( .A(n17195), .B(n23778), .X(n17193) );
  o32ai_1 U16532 ( .A1(n12505), .A2(n16979), .A3(n17196), .B1(n16974), .B2(
        n17197), .Y(n10182) );
  xnor2_1 U16533 ( .A(n17198), .B(n17199), .Y(n17197) );
  xor2_1 U16534 ( .A(n17200), .B(n23780), .X(n17199) );
  xor2_1 U16535 ( .A(n17201), .B(n17202), .X(n17196) );
  inv_1 U16536 ( .A(inData[22]), .Y(n12505) );
  o22ai_1 U16537 ( .A1(n16979), .A2(n17203), .B1(n16974), .B2(n17204), .Y(
        n10181) );
  xnor2_1 U16538 ( .A(n17205), .B(n17206), .Y(n17204) );
  xor2_1 U16539 ( .A(n23781), .B(n17207), .X(n17206) );
  inv_1 U16540 ( .A(n17208), .Y(n16974) );
  o211ai_1 U16541 ( .A1(n17209), .A2(n17210), .B1(n17119), .C1(n16677), .Y(
        n17208) );
  inv_1 U16542 ( .A(n11045), .Y(n16677) );
  a21oi_1 U16543 ( .A1(n17211), .A2(n24056), .B1(n15849), .Y(n17210) );
  inv_1 U16544 ( .A(n23679), .Y(n17203) );
  o22ai_1 U16545 ( .A1(n17212), .A2(n12660), .B1(n12663), .B2(n17213), .Y(
        n10180) );
  xor2_1 U16546 ( .A(n17214), .B(n17215), .X(n17213) );
  o21ai_0 U16547 ( .A1(n23696), .A2(n17216), .B1(n17217), .Y(n17214) );
  o32ai_1 U16548 ( .A1(n12660), .A2(n17218), .A3(n11107), .B1(n12663), .B2(
        n17219), .Y(n10179) );
  xnor2_1 U16549 ( .A(n17220), .B(n17221), .Y(n17219) );
  xor2_1 U16550 ( .A(n23691), .B(n17222), .X(n17221) );
  inv_1 U16551 ( .A(inData[10]), .Y(n11107) );
  a21oi_1 U16552 ( .A1(n17201), .A2(n23790), .B1(n17223), .Y(n17218) );
  a21oi_1 U16553 ( .A1(n23790), .A2(n23791), .B1(n17224), .Y(n17223) );
  inv_1 U16554 ( .A(n13), .Y(n17224) );
  nor2_1 U16555 ( .A(n17212), .B(n13), .Y(n17201) );
  nand2_1 U16556 ( .A(n12663), .B(n11045), .Y(n12660) );
  nand2_1 U16557 ( .A(n11084), .B(n17225), .Y(n11045) );
  o21ai_0 U16558 ( .A1(n15754), .A2(n15806), .B1(n10613), .Y(n17225) );
  inv_1 U16559 ( .A(n16680), .Y(n15806) );
  inv_1 U16560 ( .A(n15865), .Y(n15754) );
  nand2_1 U16561 ( .A(n17226), .B(n15874), .Y(n15865) );
  o211ai_1 U16562 ( .A1(n24056), .A2(n16680), .B1(n15827), .C1(n11074), .Y(
        n12663) );
  inv_1 U16563 ( .A(n17074), .Y(n11074) );
  nand3_1 U16564 ( .A(n11084), .B(n17227), .C(n17118), .Y(n17074) );
  nand2_1 U16565 ( .A(n17209), .B(n17226), .Y(n17118) );
  inv_1 U16566 ( .A(n17228), .Y(n17227) );
  nand2_1 U16567 ( .A(n17211), .B(n24058), .Y(n16680) );
  nor2_1 U16568 ( .A(n10774), .B(n17229), .Y(n10178) );
  xor2_1 U16569 ( .A(n17230), .B(n17231), .X(n17229) );
  xor2_1 U16570 ( .A(n17232), .B(n17233), .X(n17231) );
  nor2_1 U16571 ( .A(n17234), .B(n17235), .Y(n17230) );
  nand2_1 U16572 ( .A(n17236), .B(n23922), .Y(n10177) );
  xor2_1 U16573 ( .A(n17237), .B(n17238), .X(n17236) );
  mux2_1 U16574 ( .A0(n17239), .A1(n17240), .S(n17241), .X(n17238) );
  or2_0 U16575 ( .A(n45), .B(n11558), .X(n10176) );
  nand2_1 U16576 ( .A(n16206), .B(n11211), .Y(n11558) );
  o32ai_1 U16577 ( .A1(n11134), .A2(n17242), .A3(n11094), .B1(n17243), .B2(
        n11097), .Y(n10175) );
  xnor2_1 U16578 ( .A(n17244), .B(n17245), .Y(n17243) );
  o21ai_0 U16579 ( .A1(n17246), .A2(n17247), .B1(n17248), .Y(n17244) );
  xor2_1 U16580 ( .A(n23995), .B(n17249), .X(n17248) );
  nand2_1 U16581 ( .A(n11097), .B(n12681), .Y(n11094) );
  nand3_1 U16582 ( .A(n11084), .B(n15801), .C(n11360), .Y(n11097) );
  nand2_1 U16583 ( .A(n17211), .B(n15874), .Y(n15801) );
  xor2_1 U16584 ( .A(n17250), .B(n23814), .X(n17242) );
  nand2_1 U16585 ( .A(n23858), .B(n10628), .Y(n17250) );
  inv_1 U16586 ( .A(inData[30]), .Y(n11134) );
  nand2_1 U16587 ( .A(n17251), .B(n12853), .Y(n10174) );
  mux2i_1 U16588 ( .A0(n12880), .A1(n17252), .S(n12856), .Y(n17251) );
  xor2_1 U16589 ( .A(n17253), .B(n17254), .X(n17252) );
  o21ai_0 U16590 ( .A1(n17255), .A2(n17256), .B1(n17257), .Y(n17254) );
  o32ai_1 U16591 ( .A1(n17258), .A2(n11368), .A3(n10831), .B1(n11370), .B2(
        n17259), .Y(n10173) );
  xnor2_1 U16592 ( .A(n17260), .B(n17261), .Y(n17259) );
  xor2_1 U16593 ( .A(n17262), .B(n17263), .X(n17261) );
  inv_1 U16594 ( .A(inData[20]), .Y(n10831) );
  xor2_1 U16595 ( .A(n23809), .B(n23808), .X(n17258) );
  nand2_1 U16596 ( .A(n17264), .B(n12853), .Y(n10172) );
  or2_0 U16597 ( .A(n17265), .B(n12856), .X(n12853) );
  mux2i_1 U16598 ( .A0(n17266), .A1(n17267), .S(n12856), .Y(n17264) );
  inv_1 U16599 ( .A(n12863), .Y(n12856) );
  xor2_1 U16600 ( .A(n17268), .B(n17269), .X(n17267) );
  o21ai_0 U16601 ( .A1(n17270), .A2(n17271), .B1(n17272), .Y(n17268) );
  xor2_1 U16602 ( .A(n17273), .B(n12482), .X(n17266) );
  o32ai_1 U16603 ( .A1(n17274), .A2(n12866), .A3(n15898), .B1(n17275), .B2(
        n12863), .Y(n10171) );
  a21oi_1 U16604 ( .A1(n17276), .A2(n17277), .B1(n17278), .Y(n17275) );
  a21oi_1 U16605 ( .A1(n17277), .A2(n17279), .B1(n17280), .Y(n17278) );
  inv_1 U16606 ( .A(n17281), .Y(n17276) );
  inv_1 U16607 ( .A(inData[18]), .Y(n15898) );
  nand2_1 U16608 ( .A(n17265), .B(n12863), .Y(n12866) );
  nand4_1 U16609 ( .A(n17016), .B(n17282), .C(n11310), .D(n11451), .Y(n12863)
         );
  nand3_1 U16610 ( .A(n15867), .B(n24053), .C(n17283), .Y(n11451) );
  nand3_1 U16611 ( .A(n11315), .B(n24061), .C(n17011), .Y(n11310) );
  nand2_1 U16612 ( .A(n17283), .B(n17284), .Y(n17282) );
  a221oi_1 U16613 ( .A1(n11314), .A2(n17285), .B1(n17286), .B2(n15751), .C1(
        n11438), .Y(n17016) );
  nand2_1 U16614 ( .A(n17008), .B(n11308), .Y(n17265) );
  a21oi_1 U16615 ( .A1(n17286), .A2(n11438), .B1(n17284), .Y(n11308) );
  xor2_1 U16616 ( .A(n17287), .B(n17273), .X(n17274) );
  nand2_1 U16617 ( .A(n23808), .B(n17288), .Y(n17273) );
  mux2i_1 U16618 ( .A0(n17289), .A1(n17290), .S(n11360), .Y(n10170) );
  xor2_1 U16619 ( .A(n17291), .B(n17292), .X(n17290) );
  nor2_1 U16620 ( .A(n11368), .B(n17293), .Y(n17289) );
  o22ai_1 U16621 ( .A1(n11370), .A2(n17294), .B1(n11368), .B2(n17295), .Y(
        n10169) );
  xor2_1 U16622 ( .A(n17296), .B(n17297), .X(n17295) );
  xor2_1 U16623 ( .A(n17298), .B(n17299), .X(n17294) );
  or2_0 U16624 ( .A(n17300), .B(n17301), .X(n17299) );
  mux2i_1 U16625 ( .A0(n17302), .A1(n17303), .S(n11360), .Y(n10168) );
  inv_1 U16626 ( .A(n11370), .Y(n11360) );
  nand3_1 U16627 ( .A(n17304), .B(n15827), .C(n16979), .Y(n11370) );
  a21oi_1 U16628 ( .A1(n24056), .A2(n15745), .B1(n17228), .Y(n16979) );
  xor2_1 U16629 ( .A(n17305), .B(n17306), .X(n17303) );
  xor2_1 U16630 ( .A(n17307), .B(n17308), .X(n17306) );
  xor2_1 U16631 ( .A(n17309), .B(n17310), .X(n17305) );
  nor2_1 U16632 ( .A(n17311), .B(n11366), .Y(n17302) );
  or2_0 U16633 ( .A(n11355), .B(n11368), .X(n11366) );
  nor2_1 U16634 ( .A(n17312), .B(n17228), .Y(n11368) );
  nor2_1 U16635 ( .A(n15827), .B(n24056), .Y(n17228) );
  inv_1 U16636 ( .A(inData[6]), .Y(n11355) );
  xor2_1 U16637 ( .A(n17297), .B(n12478), .X(n17311) );
  nand2_1 U16638 ( .A(n755), .B(n23811), .Y(n17297) );
  o211ai_1 U16639 ( .A1(n17313), .A2(n17314), .B1(n11377), .C1(n17315), .Y(
        n10167) );
  mux2i_1 U16640 ( .A0(n17316), .A1(n17317), .S(n12442), .Y(n17315) );
  nor2_1 U16641 ( .A(n11382), .B(n17318), .Y(n17317) );
  inv_1 U16642 ( .A(n11378), .Y(n17316) );
  xor2_1 U16643 ( .A(n17319), .B(n16948), .X(n17313) );
  xor2_1 U16644 ( .A(n17320), .B(n12), .X(n17319) );
  o211ai_1 U16645 ( .A1(n12581), .A2(n11378), .B1(n11377), .C1(n17321), .Y(
        n10166) );
  mux2i_1 U16646 ( .A0(n17322), .A1(n17323), .S(n11382), .Y(n17321) );
  xor2_1 U16647 ( .A(n17324), .B(n17325), .X(n17323) );
  xor2_1 U16648 ( .A(n16583), .B(n23811), .X(n17325) );
  o21ai_0 U16649 ( .A1(n17318), .A2(n17326), .B1(inData[0]), .Y(n17322) );
  nand2_1 U16650 ( .A(n17318), .B(n17314), .Y(n11378) );
  nor2_1 U16651 ( .A(n23826), .B(n12582), .Y(n17318) );
  nand2_1 U16652 ( .A(n17327), .B(n11377), .Y(n10165) );
  or2_0 U16653 ( .A(n12717), .B(n11382), .X(n11377) );
  nand3_1 U16654 ( .A(n17328), .B(n11436), .C(n17329), .Y(n12717) );
  nor3_1 U16655 ( .A(n17285), .B(n17330), .C(n17284), .Y(n17329) );
  nand2_1 U16656 ( .A(n11453), .B(n24057), .Y(n11436) );
  inv_1 U16657 ( .A(n17331), .Y(n17328) );
  mux2i_1 U16658 ( .A0(n23826), .A1(n17332), .S(n11382), .Y(n17327) );
  inv_1 U16659 ( .A(n17314), .Y(n11382) );
  o211ai_1 U16660 ( .A1(n24059), .A2(n17333), .B1(n17334), .C1(n17335), .Y(
        n17314) );
  mux2i_1 U16661 ( .A0(n17285), .A1(n17330), .S(n15867), .Y(n17335) );
  mux2i_1 U16662 ( .A0(n17283), .A1(n15798), .S(n11314), .Y(n17334) );
  xor2_1 U16663 ( .A(n17336), .B(n17337), .X(n17332) );
  xor2_1 U16664 ( .A(n17338), .B(n17339), .X(n17337) );
  xor2_1 U16665 ( .A(n755), .B(n17340), .X(n17339) );
  xor2_1 U16666 ( .A(n17341), .B(n16507), .X(n17336) );
  o22ai_1 U16667 ( .A1(n17342), .A2(n12897), .B1(n12895), .B2(n17343), .Y(
        n10164) );
  xnor2_1 U16668 ( .A(n2116), .B(n17344), .Y(n17343) );
  nand2_1 U16669 ( .A(n23676), .B(n23702), .Y(n17344) );
  xor2_1 U16670 ( .A(n17345), .B(n16561), .X(n17342) );
  xor2_1 U16671 ( .A(n17346), .B(n12482), .X(n17345) );
  o22ai_1 U16672 ( .A1(n12897), .A2(n17347), .B1(n17348), .B2(n12895), .Y(
        n10163) );
  xor2_1 U16673 ( .A(n17349), .B(n23676), .X(n17348) );
  nand2_1 U16674 ( .A(n2116), .B(n23702), .Y(n17349) );
  xor2_1 U16675 ( .A(n17350), .B(n17351), .X(n17347) );
  xor2_1 U16676 ( .A(n17352), .B(n16516), .X(n17351) );
  xor2_1 U16677 ( .A(n17287), .B(n11668), .X(n17350) );
  o22ai_1 U16678 ( .A1(n2113), .A2(n12895), .B1(n17353), .B2(n12897), .Y(
        n10162) );
  xor2_1 U16679 ( .A(n17354), .B(n17355), .X(n17353) );
  xor2_1 U16680 ( .A(n23808), .B(n16906), .X(n17355) );
  o32ai_1 U16681 ( .A1(n12895), .A2(n17356), .A3(n11175), .B1(n12897), .B2(
        n17357), .Y(n10161) );
  xor2_1 U16682 ( .A(n17358), .B(n17359), .X(n17357) );
  xor2_1 U16683 ( .A(n17360), .B(n16550), .X(n17359) );
  xor2_1 U16684 ( .A(n17288), .B(n16742), .X(n17358) );
  inv_1 U16685 ( .A(n17361), .Y(n12897) );
  inv_1 U16686 ( .A(inData[28]), .Y(n11175) );
  o221ai_1 U16687 ( .A1(n11442), .A2(n11443), .B1(n17286), .B2(n12915), .C1(
        n17362), .Y(n12895) );
  a221oi_1 U16688 ( .A1(n17363), .A2(n24053), .B1(n17364), .B2(n15871), .C1(
        n17361), .Y(n17362) );
  nor3_1 U16689 ( .A(n11316), .B(n17331), .C(n17365), .Y(n17361) );
  o32ai_1 U16690 ( .A1(n17366), .A2(n24053), .A3(n11441), .B1(n15867), .B2(
        n11318), .Y(n17365) );
  o21ai_0 U16691 ( .A1(n11444), .A2(n11309), .B1(n17367), .Y(n17331) );
  nand3_1 U16692 ( .A(n17368), .B(n15860), .C(n12912), .Y(n11316) );
  nand2_1 U16693 ( .A(n11438), .B(n10618), .Y(n12912) );
  inv_1 U16694 ( .A(n17369), .Y(n11438) );
  nand2_1 U16695 ( .A(n17284), .B(n15871), .Y(n15860) );
  nor2_1 U16696 ( .A(n11443), .B(n24053), .Y(n17284) );
  o21ai_0 U16697 ( .A1(n15835), .A2(n11453), .B1(n17283), .Y(n17368) );
  inv_1 U16698 ( .A(n17333), .Y(n11453) );
  nand2_1 U16699 ( .A(n15856), .B(n11444), .Y(n17333) );
  inv_1 U16700 ( .A(n24053), .Y(n11444) );
  inv_1 U16701 ( .A(n11443), .Y(n15835) );
  mux2i_1 U16702 ( .A0(n11441), .A1(n24061), .S(n24059), .Y(n17364) );
  o22ai_1 U16703 ( .A1(n23860), .A2(n11226), .B1(n11617), .B2(n17370), .Y(
        n10160) );
  xnor2_1 U16704 ( .A(n17371), .B(n17372), .Y(n17370) );
  a21oi_1 U16705 ( .A1(n17373), .A2(n17374), .B1(n17375), .Y(n17371) );
  nand2_1 U16706 ( .A(n17376), .B(n12836), .Y(n10159) );
  nand2_1 U16707 ( .A(n11617), .B(n11226), .Y(n12836) );
  mux2i_1 U16708 ( .A0(n17377), .A1(n17378), .S(n11617), .Y(n17376) );
  nand3_1 U16709 ( .A(n11226), .B(n11703), .C(n11500), .Y(n11617) );
  nand2_1 U16710 ( .A(n12548), .B(n24052), .Y(n11500) );
  inv_1 U16711 ( .A(n15795), .Y(n12548) );
  xor2_1 U16712 ( .A(n23860), .B(n12510), .X(n17378) );
  xnor2_1 U16713 ( .A(n17379), .B(n17380), .Y(n17377) );
  o21ai_0 U16714 ( .A1(n17381), .A2(n17382), .B1(n17383), .Y(n17380) );
  xor2_1 U16715 ( .A(n17384), .B(n17385), .X(n17379) );
  o32ai_1 U16716 ( .A1(n11545), .A2(n17386), .A3(n11084), .B1(n11087), .B2(
        n17387), .Y(n10158) );
  xor2_1 U16717 ( .A(n17388), .B(n17389), .X(n17387) );
  xor2_1 U16718 ( .A(n17390), .B(n17391), .X(n17389) );
  nand2_1 U16719 ( .A(n17392), .B(n17393), .Y(n17390) );
  inv_1 U16720 ( .A(n17394), .Y(n17393) );
  o211ai_1 U16721 ( .A1(n10613), .A2(n15827), .B1(n17119), .C1(n12698), .Y(
        n11087) );
  inv_1 U16722 ( .A(n12681), .Y(n12698) );
  nand3_1 U16723 ( .A(n11084), .B(n16681), .C(n17304), .Y(n12681) );
  inv_1 U16724 ( .A(n17312), .Y(n17304) );
  o21ai_0 U16725 ( .A1(n24056), .A2(n17077), .B1(n17116), .Y(n17312) );
  nand2_1 U16726 ( .A(n17209), .B(n17211), .Y(n17116) );
  nor2_1 U16727 ( .A(n17395), .B(n12558), .Y(n17211) );
  inv_1 U16728 ( .A(n38), .Y(n17395) );
  nand3_1 U16729 ( .A(n12558), .B(n15874), .C(n38), .Y(n17077) );
  inv_1 U16730 ( .A(n24058), .Y(n15874) );
  nand3_1 U16731 ( .A(n38), .B(n12558), .C(n17209), .Y(n16681) );
  nand2_1 U16732 ( .A(n15745), .B(n10613), .Y(n17119) );
  inv_1 U16733 ( .A(n15740), .Y(n15745) );
  nand3_1 U16734 ( .A(n12558), .B(n24058), .C(n38), .Y(n15740) );
  nand2_1 U16735 ( .A(n24058), .B(n17226), .Y(n15827) );
  nor2_1 U16736 ( .A(n38), .B(n12558), .Y(n17226) );
  nand2_1 U16737 ( .A(n17209), .B(n15849), .Y(n11084) );
  nor2_1 U16738 ( .A(n17396), .B(n38), .Y(n15849) );
  inv_1 U16739 ( .A(n12558), .Y(n17396) );
  nor2_1 U16740 ( .A(n10613), .B(n24058), .Y(n17209) );
  inv_1 U16741 ( .A(inData[26]), .Y(n11545) );
  nand2_1 U16742 ( .A(n17397), .B(n11114), .Y(n10157) );
  nand2_1 U16743 ( .A(n11133), .B(n11117), .Y(n11114) );
  inv_1 U16744 ( .A(n15716), .Y(n11133) );
  nor2_1 U16745 ( .A(n10832), .B(n15863), .Y(n15716) );
  mux2i_1 U16746 ( .A0(n17398), .A1(n17399), .S(n11117), .Y(n17397) );
  nand2_1 U16747 ( .A(n11593), .B(n15795), .Y(n11117) );
  nand2_1 U16748 ( .A(n24062), .B(n24055), .Y(n15795) );
  nand2_1 U16749 ( .A(inData[6]), .B(n20748), .Y(n17399) );
  xor2_1 U16750 ( .A(n17400), .B(n17401), .X(n17398) );
  xor2_1 U16751 ( .A(n17402), .B(n16940), .X(n17401) );
  xor2_1 U16752 ( .A(n10627), .B(n17403), .X(n17400) );
  o21ai_0 U16753 ( .A1(n23863), .A2(n17404), .B1(n17405), .Y(n10156) );
  mux2i_1 U16754 ( .A0(n17406), .A1(n17407), .S(n12721), .Y(n17405) );
  o21ai_0 U16755 ( .A1(n2122), .A2(n17408), .B1(n17409), .Y(n17407) );
  xor2_1 U16756 ( .A(n17410), .B(n17411), .X(n17406) );
  nand2_1 U16757 ( .A(n17412), .B(n17413), .Y(n17410) );
  inv_1 U16758 ( .A(n17414), .Y(n17413) );
  o22ai_1 U16759 ( .A1(n23863), .A2(n12719), .B1(n17415), .B2(n12721), .Y(
        n10155) );
  xnor2_1 U16760 ( .A(n17416), .B(n13022), .Y(n17415) );
  o22ai_1 U16761 ( .A1(n17417), .A2(n17418), .B1(n17419), .B2(n17420), .Y(
        n13022) );
  and2_0 U16762 ( .A(n17417), .B(n17418), .X(n17419) );
  nand2_1 U16763 ( .A(n17421), .B(n13023), .Y(n17416) );
  nand2_1 U16764 ( .A(n17422), .B(n17423), .Y(n13023) );
  inv_1 U16765 ( .A(n13021), .Y(n17421) );
  xor2_1 U16766 ( .A(n12924), .B(n17424), .X(n13021) );
  nor2_1 U16767 ( .A(n17422), .B(n17423), .Y(n17424) );
  xnor2_1 U16768 ( .A(n11089), .B(n17425), .Y(n17423) );
  nor2_1 U16769 ( .A(n13024), .B(n17426), .Y(n17425) );
  inv_1 U16770 ( .A(n13025), .Y(n17426) );
  nand2_1 U16771 ( .A(n23786), .B(n17427), .Y(n13025) );
  nor2_1 U16772 ( .A(n17427), .B(n23786), .Y(n13024) );
  nor2_1 U16773 ( .A(n17428), .B(n13027), .Y(n17427) );
  nor2_1 U16774 ( .A(n17429), .B(outData[27]), .Y(n13027) );
  mux2_1 U16775 ( .A0(n11336), .A1(n17430), .S(outData[27]), .X(n17428) );
  xor2_1 U16776 ( .A(n11336), .B(n17429), .X(n17430) );
  xor2_1 U16777 ( .A(n17431), .B(n11612), .X(n17422) );
  inv_1 U16778 ( .A(n10893), .Y(n11612) );
  o22ai_1 U16779 ( .A1(n17432), .A2(n17138), .B1(n17433), .B2(n17434), .Y(
        n17431) );
  and2_0 U16780 ( .A(n17138), .B(n17432), .X(n17433) );
  inv_1 U16781 ( .A(n17435), .Y(n17432) );
  nand2_1 U16782 ( .A(n17436), .B(n12721), .Y(n12719) );
  nand2_1 U16783 ( .A(n17437), .B(n17404), .Y(n10154) );
  nand3_1 U16784 ( .A(n2122), .B(n12721), .C(n12372), .Y(n17404) );
  mux2i_1 U16785 ( .A0(n17438), .A1(n17439), .S(n12721), .Y(n17437) );
  nand2_1 U16786 ( .A(n17409), .B(inData[14]), .Y(n17439) );
  inv_1 U16787 ( .A(n17440), .Y(n17409) );
  o21ai_0 U16788 ( .A1(n2122), .A2(n12372), .B1(n17436), .Y(n17440) );
  inv_1 U16789 ( .A(n17441), .Y(n17436) );
  xnor2_1 U16790 ( .A(n17420), .B(n17442), .Y(n17438) );
  xor2_1 U16791 ( .A(n17418), .B(n17417), .X(n17442) );
  o21ai_0 U16792 ( .A1(n17443), .A2(n10625), .B1(n17444), .Y(n17417) );
  xor2_1 U16793 ( .A(n11525), .B(n17445), .X(n17444) );
  nor2_1 U16794 ( .A(n17146), .B(n17446), .Y(n17445) );
  xor2_1 U16795 ( .A(n23995), .B(n17447), .X(n17443) );
  nand2_1 U16796 ( .A(n17448), .B(n12872), .Y(n17418) );
  o211ai_1 U16797 ( .A1(n17449), .A2(n17150), .B1(n17450), .C1(n17451), .Y(
        n12872) );
  xor2_1 U16798 ( .A(n10625), .B(n17452), .X(n17451) );
  o21ai_0 U16799 ( .A1(n17453), .A2(n17454), .B1(n17142), .Y(n17450) );
  inv_1 U16800 ( .A(n23796), .Y(n17142) );
  xor2_1 U16801 ( .A(n17455), .B(n17456), .X(n17448) );
  nand2_1 U16802 ( .A(n12871), .B(n12869), .Y(n17456) );
  o21ai_0 U16803 ( .A1(n17256), .A2(n17255), .B1(n17457), .Y(n12869) );
  xor2_1 U16804 ( .A(n17458), .B(n17459), .X(n17457) );
  nand2_1 U16805 ( .A(n17257), .B(n17253), .Y(n17459) );
  o22ai_1 U16806 ( .A1(n16987), .A2(n16990), .B1(n17460), .B2(n16989), .Y(
        n17253) );
  o22ai_1 U16807 ( .A1(n12857), .A2(n12860), .B1(n17461), .B2(n12859), .Y(
        n16989) );
  o21ai_0 U16808 ( .A1(n17270), .A2(n17271), .B1(n17462), .Y(n12859) );
  xor2_1 U16809 ( .A(n17463), .B(n17464), .X(n17462) );
  and2_0 U16810 ( .A(n17272), .B(n17269), .X(n17464) );
  xor2_1 U16811 ( .A(n17465), .B(n11510), .X(n17269) );
  nand2_1 U16812 ( .A(n17277), .B(n17281), .Y(n17465) );
  nand2_1 U16813 ( .A(n17280), .B(n17279), .Y(n17281) );
  o211ai_1 U16814 ( .A1(n17466), .A2(n17467), .B1(n17468), .C1(n17469), .Y(
        n17279) );
  nand2_1 U16815 ( .A(n17470), .B(n17471), .Y(n17280) );
  o21ai_0 U16816 ( .A1(n17472), .A2(n17473), .B1(n17292), .Y(n17471) );
  xor2_1 U16817 ( .A(n17474), .B(n17475), .X(n17292) );
  o22ai_1 U16818 ( .A1(n17260), .A2(n17263), .B1(n17476), .B2(n17477), .Y(
        n17474) );
  and2_0 U16819 ( .A(n17263), .B(n17260), .X(n17477) );
  inv_1 U16820 ( .A(n17262), .Y(n17476) );
  o21ai_0 U16821 ( .A1(n17307), .A2(n17309), .B1(n17478), .Y(n17262) );
  xor2_1 U16822 ( .A(n17479), .B(n17480), .X(n17478) );
  a21oi_1 U16823 ( .A1(n17307), .A2(n17309), .B1(n17308), .Y(n17480) );
  a21oi_1 U16824 ( .A1(n17298), .A2(n17481), .B1(n17301), .Y(n17308) );
  xnor2_1 U16825 ( .A(n17482), .B(n14685), .Y(n17301) );
  nand2_1 U16826 ( .A(n17483), .B(n17484), .Y(n17482) );
  inv_1 U16827 ( .A(n17300), .Y(n17481) );
  o21ai_0 U16828 ( .A1(n17483), .A2(n17484), .B1(n24045), .Y(n17300) );
  o22ai_1 U16829 ( .A1(n17220), .A2(n17485), .B1(n17486), .B2(n17202), .Y(
        n17484) );
  inv_1 U16830 ( .A(n23790), .Y(n17202) );
  and2_0 U16831 ( .A(n17485), .B(n17220), .X(n17486) );
  mux2i_1 U16832 ( .A0(n17487), .A1(n17488), .S(n13), .Y(n17483) );
  xor2_1 U16833 ( .A(n17489), .B(n17216), .X(n17488) );
  o21ai_0 U16834 ( .A1(n17489), .A2(n17216), .B1(n17490), .Y(n17487) );
  nand2_1 U16835 ( .A(n17491), .B(n11364), .Y(n17298) );
  o211ai_1 U16836 ( .A1(n17492), .A2(n17493), .B1(n17494), .C1(n17495), .Y(
        n11364) );
  inv_1 U16837 ( .A(n17496), .Y(n17495) );
  o21ai_0 U16838 ( .A1(n12665), .A2(n17497), .B1(n10641), .Y(n17494) );
  xor2_1 U16839 ( .A(n11520), .B(n17498), .X(n17491) );
  nand2_1 U16840 ( .A(n11363), .B(n11362), .Y(n17498) );
  o21ai_0 U16841 ( .A1(n11374), .A2(n11376), .B1(n17499), .Y(n11362) );
  xor2_1 U16842 ( .A(n10936), .B(n17500), .X(n17499) );
  a21oi_1 U16843 ( .A1(n11374), .A2(n11376), .B1(n11375), .Y(n17500) );
  o22ai_1 U16844 ( .A1(n12691), .A2(n12694), .B1(n17501), .B2(n12693), .Y(
        n11375) );
  o22ai_1 U16845 ( .A1(n17502), .A2(n17503), .B1(n23714), .B2(n17504), .Y(
        n12693) );
  nor2_1 U16846 ( .A(n16705), .B(n17505), .Y(n17504) );
  xor2_1 U16847 ( .A(n17502), .B(n17506), .X(n17505) );
  and2_0 U16848 ( .A(n12694), .B(n12691), .X(n17501) );
  o22ai_1 U16849 ( .A1(n17246), .A2(n17247), .B1(n17249), .B2(n17245), .Y(
        n12694) );
  o22ai_1 U16850 ( .A1(n12684), .A2(n12687), .B1(n17507), .B2(n12685), .Y(
        n17245) );
  mux2i_1 U16851 ( .A0(n17508), .A1(n17509), .S(n23851), .Y(n12685) );
  xor2_1 U16852 ( .A(n17510), .B(n11590), .X(n17509) );
  a21oi_1 U16853 ( .A1(n11590), .A2(n17511), .B1(n17512), .Y(n17508) );
  and2_0 U16854 ( .A(n12687), .B(n12684), .X(n17507) );
  o21ai_0 U16855 ( .A1(n17513), .A2(n17514), .B1(n17515), .Y(n12687) );
  xor2_1 U16856 ( .A(n17506), .B(n17516), .X(n17513) );
  mux2_1 U16857 ( .A0(n17517), .A1(n17518), .S(n14685), .X(n12684) );
  nand2_1 U16858 ( .A(n12701), .B(n12700), .Y(n17518) );
  inv_1 U16859 ( .A(n17519), .Y(n12700) );
  xor2_1 U16860 ( .A(n17520), .B(n17521), .X(n12701) );
  o22ai_1 U16861 ( .A1(n17519), .A2(n17521), .B1(n17522), .B2(n17520), .Y(
        n17517) );
  xnor2_1 U16862 ( .A(n17523), .B(n17524), .Y(n17520) );
  xor2_1 U16863 ( .A(n17514), .B(n17525), .X(n17524) );
  inv_1 U16864 ( .A(n23856), .Y(n17514) );
  nand2_1 U16865 ( .A(n17515), .B(n17516), .Y(n17523) );
  nand2_1 U16866 ( .A(n12676), .B(n17526), .Y(n17516) );
  o21ai_0 U16867 ( .A1(n17527), .A2(n12402), .B1(n17528), .Y(n17526) );
  o211ai_1 U16868 ( .A1(n12402), .A2(n17527), .B1(n17528), .C1(n17529), .Y(
        n17515) );
  and2_0 U16869 ( .A(n17521), .B(n17519), .X(n17522) );
  o22ai_1 U16870 ( .A1(n16719), .A2(n17530), .B1(n12518), .B2(n17531), .Y(
        n17521) );
  and2_0 U16871 ( .A(n16719), .B(n17530), .X(n17531) );
  a22oi_1 U16872 ( .A1(n12829), .A2(n12832), .B1(n12831), .B2(n17532), .Y(
        n17519) );
  or2_0 U16873 ( .A(n12832), .B(n12829), .X(n17532) );
  o21ai_0 U16874 ( .A1(n12839), .A2(n17533), .B1(n17534), .Y(n12831) );
  mux2i_1 U16875 ( .A0(n12840), .A1(n17535), .S(n11570), .Y(n17533) );
  nand2_1 U16876 ( .A(n17535), .B(n17534), .Y(n12840) );
  nand2_1 U16877 ( .A(n17536), .B(n17537), .Y(n17534) );
  xor2_1 U16878 ( .A(n17538), .B(n17310), .X(n17535) );
  nor2_1 U16879 ( .A(n17537), .B(n17536), .Y(n17538) );
  xor2_1 U16880 ( .A(n17539), .B(n17540), .X(n17536) );
  xor2_1 U16881 ( .A(n23854), .B(n10942), .X(n17540) );
  o21ai_0 U16882 ( .A1(n17541), .A2(n17542), .B1(n17543), .Y(n17539) );
  xnor2_1 U16883 ( .A(n17544), .B(n16737), .Y(n17537) );
  o22ai_1 U16884 ( .A1(n16698), .A2(n17545), .B1(n23853), .B2(n17546), .Y(
        n17544) );
  nor2_1 U16885 ( .A(n17547), .B(n17548), .Y(n17546) );
  inv_1 U16886 ( .A(n17547), .Y(n17545) );
  a22oi_1 U16887 ( .A1(n17374), .A2(n17373), .B1(n17549), .B2(n17372), .Y(
        n12839) );
  xor2_1 U16888 ( .A(n17550), .B(n17551), .X(n17372) );
  a21oi_1 U16889 ( .A1(n17552), .A2(n17553), .B1(n17554), .Y(n17551) );
  a21oi_1 U16890 ( .A1(n11101), .A2(n11100), .B1(n11102), .Y(n17554) );
  o22ai_1 U16891 ( .A1(n16695), .A2(n17555), .B1(n2074), .B2(n17556), .Y(
        n11102) );
  xor2_1 U16892 ( .A(n17557), .B(n11734), .X(n17556) );
  inv_1 U16893 ( .A(n11101), .Y(n17553) );
  xor2_1 U16894 ( .A(n17558), .B(n17559), .X(n11101) );
  xor2_1 U16895 ( .A(n10630), .B(n16934), .X(n17559) );
  xor2_1 U16896 ( .A(n16716), .B(n17560), .X(n17558) );
  inv_1 U16897 ( .A(n11100), .Y(n17552) );
  nand2_1 U16898 ( .A(n17561), .B(n11112), .Y(n11100) );
  o221ai_1 U16899 ( .A1(n41), .A2(n17562), .B1(n17563), .B2(n11070), .C1(
        n17564), .Y(n11112) );
  nor2_1 U16900 ( .A(n17565), .B(n17566), .Y(n17562) );
  xnor2_1 U16901 ( .A(n16737), .B(n17567), .Y(n17561) );
  nand2_1 U16902 ( .A(n11111), .B(n11109), .Y(n17567) );
  nand2_1 U16903 ( .A(n17383), .B(n17568), .Y(n11109) );
  o21ai_0 U16904 ( .A1(n17382), .A2(n17381), .B1(n17384), .Y(n17568) );
  o21ai_0 U16905 ( .A1(n17394), .A2(n17388), .B1(n17392), .Y(n17384) );
  xor2_1 U16906 ( .A(n17391), .B(n17569), .X(n17392) );
  and2_0 U16907 ( .A(n17570), .B(n16723), .X(n17569) );
  xor2_1 U16908 ( .A(n17571), .B(n23880), .X(n17570) );
  nand4_1 U16909 ( .A(n16687), .B(n10775), .C(n10608), .D(n15913), .Y(n17388)
         );
  nor2_1 U16910 ( .A(n16723), .B(n17572), .Y(n17394) );
  a21oi_1 U16911 ( .A1(n17571), .A2(n23880), .B1(n17382), .Y(n17572) );
  xnor2_1 U16912 ( .A(n17573), .B(n17574), .Y(n17383) );
  and2_0 U16913 ( .A(n17381), .B(n17382), .X(n17574) );
  nor2_1 U16914 ( .A(n17571), .B(n23880), .Y(n17382) );
  nand2_1 U16915 ( .A(n17575), .B(n17576), .Y(n17571) );
  xor2_1 U16916 ( .A(n11574), .B(n17577), .X(n17575) );
  nand2_1 U16917 ( .A(outData[3]), .B(n17578), .Y(n17577) );
  xor2_1 U16918 ( .A(n17579), .B(n17580), .X(n17381) );
  xor2_1 U16919 ( .A(n41), .B(n17563), .X(n17580) );
  xor2_1 U16920 ( .A(n16801), .B(n11070), .X(n17579) );
  o211ai_1 U16921 ( .A1(n17565), .A2(n17566), .B1(n17581), .C1(n17582), .Y(
        n11111) );
  inv_1 U16922 ( .A(n17564), .Y(n17582) );
  o21ai_0 U16923 ( .A1(n16695), .A2(n17583), .B1(n17584), .Y(n17564) );
  mux2i_1 U16924 ( .A0(n17585), .A1(n17557), .S(n17586), .Y(n17584) );
  and2_0 U16925 ( .A(n16695), .B(n17555), .X(n17557) );
  nor2_1 U16926 ( .A(n17587), .B(n17555), .Y(n17585) );
  xnor2_1 U16927 ( .A(n17555), .B(n17586), .Y(n17583) );
  xor2_1 U16928 ( .A(n17588), .B(n2074), .X(n17586) );
  xnor2_1 U16929 ( .A(n16801), .B(n17589), .Y(n17555) );
  xor2_1 U16930 ( .A(n12440), .B(n17590), .X(n17589) );
  o21ai_0 U16931 ( .A1(n17563), .A2(n11070), .B1(n41), .Y(n17581) );
  inv_1 U16932 ( .A(n17563), .Y(n17566) );
  a21oi_1 U16933 ( .A1(n17576), .A2(outData[4]), .B1(n17590), .Y(n17563) );
  inv_1 U16934 ( .A(n17375), .Y(n17549) );
  xor2_1 U16935 ( .A(n17591), .B(n17592), .X(n17375) );
  nor2_1 U16936 ( .A(n17373), .B(n17374), .Y(n17592) );
  xor2_1 U16937 ( .A(n17593), .B(n17594), .X(n17373) );
  xor2_1 U16938 ( .A(n23853), .B(n17595), .X(n17594) );
  xor2_1 U16939 ( .A(n17548), .B(n17547), .X(n17593) );
  nor2_1 U16940 ( .A(n17596), .B(n17597), .Y(n17547) );
  xnor2_1 U16941 ( .A(n17598), .B(n17599), .Y(n17596) );
  nand2_1 U16942 ( .A(outData[7]), .B(n17600), .Y(n17599) );
  o22ai_1 U16943 ( .A1(n16716), .A2(n17601), .B1(n17602), .B2(n10630), .Y(
        n17374) );
  nor2_1 U16944 ( .A(n17560), .B(n17603), .Y(n17602) );
  inv_1 U16945 ( .A(n17601), .Y(n17560) );
  o21ai_0 U16946 ( .A1(n17604), .A2(n10619), .B1(n17600), .Y(n17601) );
  and2_0 U16947 ( .A(n12440), .B(n17590), .X(n17604) );
  xor2_1 U16948 ( .A(n17605), .B(n17530), .X(n12832) );
  xor2_1 U16949 ( .A(n11520), .B(n17606), .X(n17530) );
  a21oi_1 U16950 ( .A1(n17607), .A2(outData[9]), .B1(n17527), .Y(n17606) );
  xor2_1 U16951 ( .A(n16719), .B(n12518), .X(n17605) );
  xor2_1 U16952 ( .A(n17608), .B(n11292), .X(n12829) );
  nand2_1 U16953 ( .A(n17609), .B(n17610), .Y(n17608) );
  o21ai_0 U16954 ( .A1(n17541), .A2(n17542), .B1(n23854), .Y(n17610) );
  xor2_1 U16955 ( .A(n17543), .B(n17611), .X(n17609) );
  nand2_1 U16956 ( .A(n17541), .B(n17542), .Y(n17543) );
  xor2_1 U16957 ( .A(n12330), .B(n17597), .X(n17542) );
  and2_0 U16958 ( .A(n17246), .B(n17247), .X(n17249) );
  xor2_1 U16959 ( .A(n17612), .B(n17613), .X(n17247) );
  inv_1 U16960 ( .A(n17502), .Y(n17613) );
  xnor2_1 U16961 ( .A(n17614), .B(n17615), .Y(n17502) );
  xor2_1 U16962 ( .A(n17616), .B(outData[12]), .X(n17614) );
  xor2_1 U16963 ( .A(n16705), .B(n23714), .X(n17612) );
  inv_1 U16964 ( .A(n17617), .Y(n17246) );
  o22ai_1 U16965 ( .A1(n17618), .A2(n17510), .B1(n23851), .B2(n17619), .Y(
        n17617) );
  xor2_1 U16966 ( .A(n17620), .B(n17512), .X(n17619) );
  nor2_1 U16967 ( .A(n11590), .B(n17511), .Y(n17512) );
  inv_1 U16968 ( .A(n17510), .Y(n17511) );
  inv_1 U16969 ( .A(n17618), .Y(n11590) );
  nand2_1 U16970 ( .A(n17621), .B(n17615), .Y(n17510) );
  xor2_1 U16971 ( .A(n13014), .B(n17622), .X(n17621) );
  nand2_1 U16972 ( .A(outData[11]), .B(n17528), .Y(n17622) );
  xnor2_1 U16973 ( .A(n17623), .B(n17624), .Y(n12691) );
  xor2_1 U16974 ( .A(n23789), .B(n16737), .X(n17624) );
  xor2_1 U16975 ( .A(n12671), .B(n17625), .X(n17623) );
  o22ai_1 U16976 ( .A1(n17625), .A2(n12671), .B1(n23789), .B2(n17626), .Y(
        n11376) );
  and2_0 U16977 ( .A(n12671), .B(n17625), .X(n17626) );
  a211oi_1 U16978 ( .A1(n17615), .A2(outData[13]), .B1(n17627), .C1(n11173), 
        .Y(n17625) );
  xor2_1 U16979 ( .A(n17628), .B(n17629), .X(n11374) );
  xor2_1 U16980 ( .A(n23788), .B(n12297), .X(n17629) );
  xor2_1 U16981 ( .A(n17493), .B(n17492), .X(n17628) );
  o211ai_1 U16982 ( .A1(n12665), .A2(n17497), .B1(n17630), .C1(n17496), .Y(
        n11363) );
  xnor2_1 U16983 ( .A(n17631), .B(n17220), .Y(n17496) );
  xor2_1 U16984 ( .A(n17485), .B(n23790), .X(n17631) );
  o21ai_0 U16985 ( .A1(n17632), .A2(n17633), .B1(n17634), .Y(n17485) );
  o21ai_0 U16986 ( .A1(n17492), .A2(n17493), .B1(n23788), .Y(n17630) );
  inv_1 U16987 ( .A(n17492), .Y(n17497) );
  a21oi_1 U16988 ( .A1(n17635), .A2(outData[14]), .B1(n17632), .Y(n17492) );
  xnor2_1 U16989 ( .A(n17636), .B(n17637), .Y(n17309) );
  xor2_1 U16990 ( .A(n17212), .B(n17207), .X(n17636) );
  inv_1 U16991 ( .A(n17638), .Y(n17207) );
  and2_0 U16992 ( .A(n17639), .B(n17640), .X(n17307) );
  o21ai_0 U16993 ( .A1(n17489), .A2(n17216), .B1(n13), .Y(n17640) );
  xor2_1 U16994 ( .A(n16904), .B(n17490), .X(n17639) );
  nand2_1 U16995 ( .A(n17489), .B(n17216), .Y(n17490) );
  xor2_1 U16996 ( .A(outData[16]), .B(n17634), .X(n17489) );
  xnor2_1 U16997 ( .A(n17198), .B(n17641), .Y(n17263) );
  xor2_1 U16998 ( .A(n23679), .B(n17642), .X(n17641) );
  xor2_1 U16999 ( .A(n17643), .B(n17588), .X(n17260) );
  inv_1 U17000 ( .A(n17644), .Y(n17588) );
  o22ai_1 U17001 ( .A1(n17638), .A2(n17637), .B1(n17645), .B2(n17212), .Y(
        n17643) );
  inv_1 U17002 ( .A(n23791), .Y(n17212) );
  and2_0 U17003 ( .A(n17637), .B(n17638), .X(n17645) );
  o21ai_0 U17004 ( .A1(n12346), .A2(n17646), .B1(n17647), .Y(n17637) );
  mux2i_1 U17005 ( .A0(n17648), .A1(n17649), .S(n17650), .Y(n17470) );
  o21ai_0 U17006 ( .A1(n10942), .A2(n17651), .B1(n17652), .Y(n17649) );
  xnor2_1 U17007 ( .A(n17473), .B(n17472), .Y(n17651) );
  inv_1 U17008 ( .A(n17291), .Y(n17648) );
  o211ai_1 U17009 ( .A1(n17472), .A2(n17473), .B1(n17653), .C1(n17652), .Y(
        n17291) );
  nand3_1 U17010 ( .A(n17472), .B(n17473), .C(n10942), .Y(n17652) );
  inv_1 U17011 ( .A(n17654), .Y(n17653) );
  a21oi_1 U17012 ( .A1(n17473), .A2(n17472), .B1(n10942), .Y(n17654) );
  o22ai_1 U17013 ( .A1(n17642), .A2(n17198), .B1(n23679), .B2(n17655), .Y(
        n17473) );
  and2_0 U17014 ( .A(n17198), .B(n17642), .X(n17655) );
  a21oi_1 U17015 ( .A1(n17647), .A2(outData[18]), .B1(n17656), .Y(n17642) );
  xnor2_1 U17016 ( .A(n17657), .B(n17658), .Y(n17472) );
  xor2_1 U17017 ( .A(n12544), .B(n16898), .X(n17658) );
  xor2_1 U17018 ( .A(n17467), .B(n17659), .X(n17657) );
  inv_1 U17019 ( .A(n17660), .Y(n17277) );
  a211oi_1 U17020 ( .A1(n17468), .A2(n17467), .B1(n17466), .C1(n17469), .Y(
        n17660) );
  xnor2_1 U17021 ( .A(n17661), .B(n17662), .Y(n17469) );
  xor2_1 U17022 ( .A(n16985), .B(n16707), .X(n17662) );
  nand2_1 U17023 ( .A(n17663), .B(n17664), .Y(n17661) );
  nor2_1 U17024 ( .A(n17665), .B(n12544), .Y(n17466) );
  xor2_1 U17025 ( .A(n24045), .B(n17659), .X(n17665) );
  inv_1 U17026 ( .A(n17666), .Y(n17659) );
  nand2_1 U17027 ( .A(n12544), .B(n17666), .Y(n17468) );
  o21ai_0 U17028 ( .A1(n17656), .A2(n17051), .B1(n17667), .Y(n17666) );
  nand2_1 U17029 ( .A(n17270), .B(n17271), .Y(n17272) );
  mux2i_1 U17030 ( .A0(n17668), .A1(n17669), .S(n23697), .Y(n17271) );
  o21ai_0 U17031 ( .A1(n17670), .A2(n17671), .B1(n17672), .Y(n17669) );
  xor2_1 U17032 ( .A(n17670), .B(n17671), .X(n17668) );
  a21oi_1 U17033 ( .A1(n16985), .A2(n17663), .B1(n17673), .Y(n17270) );
  inv_1 U17034 ( .A(n17664), .Y(n17673) );
  nand2_1 U17035 ( .A(n17674), .B(n16975), .Y(n17664) );
  or2_0 U17036 ( .A(n17674), .B(n16975), .X(n17663) );
  xor2_1 U17037 ( .A(n17675), .B(n17676), .X(n17674) );
  inv_1 U17038 ( .A(n23793), .Y(n16985) );
  and2_0 U17039 ( .A(n12860), .B(n12857), .X(n17461) );
  o22ai_1 U17040 ( .A1(n17670), .A2(n17671), .B1(n17677), .B2(n17678), .Y(
        n12860) );
  inv_1 U17041 ( .A(n23697), .Y(n17678) );
  xor2_1 U17042 ( .A(n17679), .B(n17672), .X(n17677) );
  nand2_1 U17043 ( .A(n17670), .B(n17671), .Y(n17672) );
  xor2_1 U17044 ( .A(n17680), .B(n17616), .X(n17671) );
  o211ai_1 U17045 ( .A1(n17675), .A2(n11468), .B1(n12977), .C1(n17681), .Y(
        n17680) );
  nand2_1 U17046 ( .A(outData[21]), .B(outData[20]), .Y(n12977) );
  xnor2_1 U17047 ( .A(n17682), .B(n17683), .Y(n12857) );
  xor2_1 U17048 ( .A(n23794), .B(n17684), .X(n17683) );
  and2_0 U17049 ( .A(n16990), .B(n16987), .X(n17460) );
  o22ai_1 U17050 ( .A1(n17684), .A2(n17682), .B1(n17685), .B2(n16983), .Y(
        n16990) );
  inv_1 U17051 ( .A(n23794), .Y(n16983) );
  and2_0 U17052 ( .A(n17682), .B(n17684), .X(n17685) );
  a21oi_1 U17053 ( .A1(outData[22]), .A2(n17681), .B1(n17686), .Y(n17684) );
  mux2_1 U17054 ( .A0(n17687), .A1(n17688), .S(n23795), .X(n16987) );
  o21ai_0 U17055 ( .A1(n17689), .A2(n17690), .B1(n17691), .Y(n17688) );
  xor2_1 U17056 ( .A(n17132), .B(n17692), .X(n17687) );
  xnor2_1 U17057 ( .A(n11668), .B(n17693), .Y(n17257) );
  and2_0 U17058 ( .A(n17255), .B(n17256), .X(n17693) );
  xnor2_1 U17059 ( .A(n17694), .B(n17454), .Y(n17255) );
  xor2_1 U17060 ( .A(n17453), .B(n23796), .X(n17694) );
  inv_1 U17061 ( .A(n17695), .Y(n17256) );
  o22ai_1 U17062 ( .A1(n17689), .A2(n17690), .B1(n23795), .B2(n17696), .Y(
        n17695) );
  xor2_1 U17063 ( .A(n17697), .B(n17691), .X(n17696) );
  nand2_1 U17064 ( .A(n17689), .B(n17690), .Y(n17691) );
  inv_1 U17065 ( .A(n17692), .Y(n17690) );
  a21oi_1 U17066 ( .A1(outData[23]), .A2(n17698), .B1(n17699), .Y(n17692) );
  xnor2_1 U17067 ( .A(n17700), .B(n11103), .Y(n12871) );
  o211ai_1 U17068 ( .A1(n17453), .A2(n17454), .B1(n17701), .C1(n17702), .Y(
        n17700) );
  xor2_1 U17069 ( .A(n17452), .B(n23766), .X(n17702) );
  o21ai_0 U17070 ( .A1(n17146), .A2(n17446), .B1(n17447), .Y(n17452) );
  nand2_1 U17071 ( .A(n17146), .B(n17446), .Y(n17447) );
  nand2_1 U17072 ( .A(n17703), .B(n17704), .Y(n17446) );
  inv_1 U17073 ( .A(n17705), .Y(n17704) );
  xor2_1 U17074 ( .A(n17133), .B(n17706), .X(n17703) );
  nand2_1 U17075 ( .A(outData[25]), .B(n17707), .Y(n17706) );
  o21ai_0 U17076 ( .A1(n17449), .A2(n17150), .B1(n23796), .Y(n17701) );
  inv_1 U17077 ( .A(n17449), .Y(n17454) );
  xnor2_1 U17078 ( .A(n17708), .B(n10796), .Y(n17449) );
  o21ai_0 U17079 ( .A1(n17699), .A2(n17709), .B1(n17707), .Y(n17708) );
  xnor2_1 U17080 ( .A(n17138), .B(n17710), .Y(n17420) );
  xor2_1 U17081 ( .A(n17434), .B(n17435), .X(n17710) );
  o21ai_0 U17082 ( .A1(n17705), .A2(n17711), .B1(n17429), .Y(n17435) );
  xnor2_1 U17083 ( .A(n17712), .B(n16898), .Y(n17429) );
  nand2_1 U17084 ( .A(n17705), .B(n17711), .Y(n17712) );
  nor2_1 U17085 ( .A(n17707), .B(outData[25]), .Y(n17705) );
  nand2_1 U17086 ( .A(n17699), .B(n17709), .Y(n17707) );
  nor2_1 U17087 ( .A(n17698), .B(outData[23]), .Y(n17699) );
  inv_1 U17088 ( .A(n17686), .Y(n17698) );
  xor2_1 U17089 ( .A(n17644), .B(n17713), .X(n17686) );
  nor2_1 U17090 ( .A(outData[22]), .B(n17681), .Y(n17713) );
  nand3_1 U17091 ( .A(n17676), .B(n11468), .C(n17675), .Y(n17681) );
  inv_1 U17092 ( .A(n17667), .Y(n17675) );
  nand2_1 U17093 ( .A(n17656), .B(n17051), .Y(n17667) );
  nor2_1 U17094 ( .A(n17647), .B(outData[18]), .Y(n17656) );
  nand2_1 U17095 ( .A(n17646), .B(n12346), .Y(n17647) );
  nor2_1 U17096 ( .A(n17634), .B(outData[16]), .Y(n17646) );
  xnor2_1 U17097 ( .A(n17714), .B(n17715), .Y(n17634) );
  nand2_1 U17098 ( .A(n17632), .B(n17633), .Y(n17714) );
  nor2_1 U17099 ( .A(n17635), .B(outData[14]), .Y(n17632) );
  inv_1 U17100 ( .A(n17627), .Y(n17635) );
  nor3_1 U17101 ( .A(outData[13]), .B(outData[12]), .C(n17615), .Y(n17627) );
  or2_0 U17102 ( .A(n17528), .B(outData[11]), .X(n17615) );
  nand2_1 U17103 ( .A(n17527), .B(n12402), .Y(n17528) );
  nor2_1 U17104 ( .A(n17607), .B(outData[9]), .Y(n17527) );
  nand2_1 U17105 ( .A(n17597), .B(n12330), .Y(n17607) );
  nor2_1 U17106 ( .A(n17600), .B(outData[7]), .Y(n17597) );
  nand3_1 U17107 ( .A(n12440), .B(n10619), .C(n17590), .Y(n17600) );
  nor2_1 U17108 ( .A(n17576), .B(outData[4]), .Y(n17590) );
  nand2_1 U17109 ( .A(n17716), .B(n12354), .Y(n17576) );
  inv_1 U17110 ( .A(n17578), .Y(n17716) );
  inv_1 U17111 ( .A(n23787), .Y(n17434) );
  mux2i_1 U17112 ( .A0(n17717), .A1(n17718), .S(n12721), .Y(n10153) );
  o221ai_1 U17113 ( .A1(n24061), .A2(n11318), .B1(n12915), .B2(n17719), .C1(
        n17369), .Y(n12721) );
  nand2_1 U17114 ( .A(n15798), .B(n11445), .Y(n17369) );
  mux2i_1 U17115 ( .A0(n15867), .A1(n20751), .S(n24053), .Y(n17719) );
  nor3_1 U17116 ( .A(n17720), .B(n17441), .C(n12699), .Y(n17718) );
  inv_1 U17117 ( .A(inData[24]), .Y(n12699) );
  a221oi_1 U17118 ( .A1(n17721), .A2(n24061), .B1(n15867), .B2(n17285), .C1(
        n17363), .Y(n17441) );
  inv_1 U17119 ( .A(n11320), .Y(n15867) );
  nand2_1 U17120 ( .A(n10618), .B(n17286), .Y(n11320) );
  nand2_1 U17121 ( .A(n15871), .B(n17011), .Y(n17721) );
  inv_1 U17122 ( .A(n11454), .Y(n17011) );
  xor2_1 U17123 ( .A(n23815), .B(n12372), .X(n17720) );
  xnor2_1 U17124 ( .A(n17722), .B(n17723), .Y(n17717) );
  o21ai_0 U17125 ( .A1(n16414), .A2(n11106), .B1(n17724), .Y(n17723) );
  o22ai_1 U17126 ( .A1(n23924), .A2(n11331), .B1(n17725), .B2(n11333), .Y(
        n10152) );
  xor2_1 U17127 ( .A(n17726), .B(n17727), .X(n17725) );
  xor2_1 U17128 ( .A(n16832), .B(n17728), .X(n17727) );
  nand2_1 U17129 ( .A(n17729), .B(n17730), .Y(n17728) );
  nand2_1 U17130 ( .A(n11333), .B(n12792), .Y(n11331) );
  nand3_1 U17131 ( .A(n11443), .B(n17367), .C(n17731), .Y(n12792) );
  inv_1 U17132 ( .A(n17732), .Y(n17731) );
  o22ai_1 U17133 ( .A1(n11309), .A2(n11454), .B1(n11311), .B2(n11319), .Y(
        n17732) );
  xnor2_1 U17134 ( .A(n10618), .B(n24053), .Y(n11454) );
  nand2_1 U17135 ( .A(n17283), .B(n17286), .Y(n11309) );
  inv_1 U17136 ( .A(n12915), .Y(n17283) );
  nand3_1 U17137 ( .A(n24061), .B(n15871), .C(n24059), .Y(n17367) );
  nand2_1 U17138 ( .A(n20751), .B(n24061), .Y(n11443) );
  o211ai_1 U17139 ( .A1(n17733), .A2(n17286), .B1(n17734), .C1(n17008), .Y(
        n11333) );
  a21oi_1 U17140 ( .A1(n15751), .A2(n15856), .B1(n17363), .Y(n17008) );
  nor2_1 U17141 ( .A(n12915), .B(n11319), .Y(n17363) );
  nand2_1 U17142 ( .A(n24057), .B(n24059), .Y(n12915) );
  inv_1 U17143 ( .A(n11319), .Y(n15856) );
  nand2_1 U17144 ( .A(n20751), .B(n17286), .Y(n11319) );
  o21ai_0 U17145 ( .A1(n15798), .A2(n17330), .B1(n11314), .Y(n17734) );
  inv_1 U17146 ( .A(n11441), .Y(n11314) );
  nand2_1 U17147 ( .A(n24061), .B(n10618), .Y(n11441) );
  inv_1 U17148 ( .A(n11311), .Y(n17330) );
  nand2_1 U17149 ( .A(n15751), .B(n11445), .Y(n11311) );
  nor2_1 U17150 ( .A(n24053), .B(n24057), .Y(n15798) );
  inv_1 U17151 ( .A(n24061), .Y(n17286) );
  a21oi_1 U17152 ( .A1(n11315), .A2(n24053), .B1(n17285), .Y(n17733) );
  inv_1 U17153 ( .A(n11318), .Y(n17285) );
  nand2_1 U17154 ( .A(n24059), .B(n15751), .Y(n11318) );
  inv_1 U17155 ( .A(n11442), .Y(n15751) );
  nand2_1 U17156 ( .A(n24053), .B(n15871), .Y(n11442) );
  inv_1 U17157 ( .A(n24057), .Y(n15871) );
  inv_1 U17158 ( .A(n17366), .Y(n11315) );
  nand2_1 U17159 ( .A(n24057), .B(n11445), .Y(n17366) );
  inv_1 U17160 ( .A(n24059), .Y(n11445) );
  nand2_1 U17161 ( .A(n23922), .B(n17735), .Y(n10151) );
  xnor2_1 U17162 ( .A(n16223), .B(n17736), .Y(n17735) );
  xor2_1 U17163 ( .A(n16224), .B(n17737), .X(n17736) );
  o22ai_1 U17164 ( .A1(n17738), .A2(n16730), .B1(n60), .B2(n17739), .Y(n16224)
         );
  nor2_1 U17165 ( .A(n11755), .B(n11757), .Y(n17739) );
  inv_1 U17166 ( .A(n11757), .Y(n17738) );
  o22ai_1 U17167 ( .A1(n13031), .A2(n13029), .B1(n23803), .B2(n17740), .Y(
        n11757) );
  and2_0 U17168 ( .A(n13029), .B(n13031), .X(n17740) );
  o22ai_1 U17169 ( .A1(n11763), .A2(n11765), .B1(n17741), .B2(n17742), .Y(
        n13029) );
  inv_1 U17170 ( .A(n23804), .Y(n17742) );
  and2_0 U17171 ( .A(n11765), .B(n11763), .X(n17741) );
  o22ai_1 U17172 ( .A1(n11631), .A2(n11632), .B1(n59), .B2(n17743), .Y(n11765)
         );
  and2_0 U17173 ( .A(n11632), .B(n11631), .X(n17743) );
  o22ai_1 U17174 ( .A1(n16872), .A2(n16996), .B1(n12372), .B2(n17744), .Y(
        n11632) );
  and2_0 U17175 ( .A(n16996), .B(n16872), .X(n17744) );
  xor2_1 U17176 ( .A(n17745), .B(n17746), .X(n16996) );
  o21ai_0 U17177 ( .A1(n23815), .A2(n16277), .B1(n17747), .Y(n17745) );
  xor2_1 U17178 ( .A(n17650), .B(n17748), .X(n17747) );
  nor2_1 U17179 ( .A(n17005), .B(n17001), .Y(n17748) );
  a21oi_1 U17180 ( .A1(n16882), .A2(n12546), .B1(n17749), .Y(n17001) );
  xor2_1 U17181 ( .A(n17591), .B(n17750), .X(n17749) );
  a21oi_1 U17182 ( .A1(n12879), .A2(n12880), .B1(n12878), .Y(n17750) );
  o22ai_1 U17183 ( .A1(n12890), .A2(n17751), .B1(n17752), .B2(n12862), .Y(
        n12878) );
  inv_1 U17184 ( .A(n10), .Y(n12862) );
  nor2_1 U17185 ( .A(n12891), .B(n16894), .Y(n17752) );
  inv_1 U17186 ( .A(n17751), .Y(n12891) );
  o21ai_0 U17187 ( .A1(n16637), .A2(n12902), .B1(n17753), .Y(n17751) );
  xor2_1 U17188 ( .A(n17479), .B(n17754), .X(n17753) );
  a21oi_1 U17189 ( .A1(n12902), .A2(n16637), .B1(n12900), .Y(n17754) );
  o22ai_1 U17190 ( .A1(n12907), .A2(n12906), .B1(n17755), .B2(n17756), .Y(
        n12900) );
  inv_1 U17191 ( .A(n9), .Y(n17756) );
  and2_0 U17192 ( .A(n12906), .B(n12907), .X(n17755) );
  xnor2_1 U17193 ( .A(n17757), .B(n17758), .Y(n12906) );
  o21ai_0 U17194 ( .A1(n6), .A2(n16516), .B1(n17759), .Y(n17757) );
  xor2_1 U17195 ( .A(n11520), .B(n17760), .X(n17759) );
  o21ai_0 U17196 ( .A1(n17287), .A2(n17761), .B1(n17352), .Y(n17760) );
  o22ai_1 U17197 ( .A1(n16906), .A2(n17762), .B1(n17763), .B2(n17293), .Y(
        n17352) );
  inv_1 U17198 ( .A(n23808), .Y(n17293) );
  nor2_1 U17199 ( .A(n16542), .B(n17354), .Y(n17763) );
  inv_1 U17200 ( .A(n17354), .Y(n17762) );
  xor2_1 U17201 ( .A(n17764), .B(n17765), .X(n17354) );
  o22ai_1 U17202 ( .A1(n17766), .A2(n17360), .B1(n17767), .B2(n17288), .Y(
        n17764) );
  inv_1 U17203 ( .A(n23809), .Y(n17288) );
  and2_0 U17204 ( .A(n17360), .B(n17766), .X(n17767) );
  o22ai_1 U17205 ( .A1(n16912), .A2(n17346), .B1(n17768), .B2(n17769), .Y(
        n17360) );
  inv_1 U17206 ( .A(n12482), .Y(n17769) );
  and2_0 U17207 ( .A(n17346), .B(n16912), .X(n17768) );
  o22ai_1 U17208 ( .A1(n16916), .A2(n17320), .B1(n17770), .B2(n17296), .Y(
        n17346) );
  inv_1 U17209 ( .A(n12), .Y(n17296) );
  and2_0 U17210 ( .A(n17320), .B(n16916), .X(n17770) );
  o22ai_1 U17211 ( .A1(n16583), .A2(n17771), .B1(n17772), .B2(n11365), .Y(
        n17320) );
  inv_1 U17212 ( .A(n23811), .Y(n11365) );
  nor2_1 U17213 ( .A(n17324), .B(n16921), .Y(n17772) );
  inv_1 U17214 ( .A(n17324), .Y(n17771) );
  xnor2_1 U17215 ( .A(n17773), .B(n17774), .Y(n17324) );
  o22ai_1 U17216 ( .A1(n17775), .A2(n16507), .B1(n755), .B2(n17776), .Y(n17773) );
  nor2_1 U17217 ( .A(n17777), .B(n17341), .Y(n17776) );
  inv_1 U17218 ( .A(n17341), .Y(n17775) );
  o22ai_1 U17219 ( .A1(n11386), .A2(n11385), .B1(n12478), .B2(n17778), .Y(
        n17341) );
  and2_0 U17220 ( .A(n11385), .B(n11386), .X(n17778) );
  o22ai_1 U17221 ( .A1(n12705), .A2(n12708), .B1(n17779), .B2(n12707), .Y(
        n11385) );
  inv_1 U17222 ( .A(n23814), .Y(n12707) );
  and2_0 U17223 ( .A(n12708), .B(n12705), .X(n17779) );
  o22ai_1 U17224 ( .A1(n17780), .A2(n12715), .B1(n23858), .B2(n17781), .Y(
        n12708) );
  nor2_1 U17225 ( .A(n12640), .B(n12716), .Y(n17781) );
  inv_1 U17226 ( .A(n12716), .Y(n17780) );
  o22ai_1 U17227 ( .A1(n16933), .A2(n11129), .B1(n17782), .B2(n10628), .Y(
        n12716) );
  and2_0 U17228 ( .A(n11129), .B(n16933), .X(n17782) );
  o21ai_0 U17229 ( .A1(n23715), .A2(n17783), .B1(n17784), .Y(n11129) );
  xor2_1 U17230 ( .A(n17031), .B(n17785), .X(n17784) );
  o21ai_0 U17231 ( .A1(n12690), .A2(n12725), .B1(n12724), .Y(n17785) );
  o22ai_1 U17232 ( .A1(n16938), .A2(n11138), .B1(n17786), .B2(n12838), .Y(
        n12724) );
  inv_1 U17233 ( .A(n23712), .Y(n12838) );
  and2_0 U17234 ( .A(n11138), .B(n16938), .X(n17786) );
  o22ai_1 U17235 ( .A1(n12443), .A2(n17402), .B1(n17787), .B2(n10627), .Y(
        n11138) );
  and2_0 U17236 ( .A(n17402), .B(n12443), .X(n17787) );
  o21ai_0 U17237 ( .A1(n16674), .A2(n17788), .B1(n17789), .Y(n17402) );
  xor2_1 U17238 ( .A(n11570), .B(n17790), .X(n17789) );
  a21oi_1 U17239 ( .A1(n16674), .A2(n17788), .B1(n12732), .Y(n17790) );
  a21oi_1 U17240 ( .A1(n16415), .A2(n12487), .B1(n17791), .Y(n12732) );
  xor2_1 U17241 ( .A(n11301), .B(n17792), .X(n17791) );
  nand2_1 U17242 ( .A(n17722), .B(n17724), .Y(n17792) );
  nand2_1 U17243 ( .A(n16414), .B(n11106), .Y(n17724) );
  inv_1 U17244 ( .A(n12487), .Y(n11106) );
  a22oi_1 U17245 ( .A1(n17793), .A2(n11122), .B1(n17386), .B2(n17794), .Y(
        n17722) );
  or2_0 U17246 ( .A(n11122), .B(n17793), .X(n17794) );
  inv_1 U17247 ( .A(n23861), .Y(n17386) );
  a21oi_1 U17248 ( .A1(n17412), .A2(n17411), .B1(n17414), .Y(n11122) );
  nor2_1 U17249 ( .A(n16391), .B(n19), .Y(n17414) );
  nor2_1 U17250 ( .A(n11105), .B(n11531), .Y(n17411) );
  inv_1 U17251 ( .A(n23687), .Y(n11105) );
  nand2_1 U17252 ( .A(n19), .B(n16391), .Y(n17412) );
  inv_1 U17253 ( .A(n12510), .Y(n17788) );
  inv_1 U17254 ( .A(n23715), .Y(n12690) );
  inv_1 U17255 ( .A(n6), .Y(n17287) );
  inv_1 U17256 ( .A(n11), .Y(n12902) );
  inv_1 U17257 ( .A(n12546), .Y(n12880) );
  nor2_1 U17258 ( .A(n17004), .B(n17003), .Y(n17005) );
  inv_1 U17259 ( .A(n23815), .Y(n17004) );
  inv_1 U17260 ( .A(n17616), .Y(n17650) );
  xor2_1 U17261 ( .A(n16228), .B(n16226), .X(n16223) );
  inv_1 U17262 ( .A(n12452), .Y(n16228) );
  nand2_1 U17263 ( .A(n11593), .B(n17795), .Y(n10150) );
  xnor2_1 U17264 ( .A(n17796), .B(n17797), .Y(n17795) );
  xnor2_1 U17265 ( .A(n17798), .B(n17799), .Y(n17797) );
  nand2_1 U17266 ( .A(n11593), .B(n17800), .Y(n10149) );
  xnor2_1 U17267 ( .A(n17801), .B(n17802), .Y(n17800) );
  xor2_1 U17268 ( .A(n17803), .B(n17804), .X(n17802) );
  nand2_1 U17269 ( .A(n11593), .B(n17805), .Y(n10148) );
  xor2_1 U17270 ( .A(n17806), .B(n17807), .X(n17805) );
  xor2_1 U17271 ( .A(n10814), .B(n17679), .X(n17807) );
  inv_1 U17272 ( .A(n17031), .Y(n17679) );
  o22ai_1 U17273 ( .A1(n17804), .A2(n17803), .B1(n17808), .B2(n17801), .Y(
        n10814) );
  xnor2_1 U17274 ( .A(n17809), .B(n13368), .Y(n17801) );
  o22ai_1 U17275 ( .A1(n16730), .A2(n17810), .B1(n17811), .B2(n17812), .Y(
        n17809) );
  inv_1 U17276 ( .A(n23875), .Y(n17812) );
  nor2_1 U17277 ( .A(n12351), .B(n11755), .Y(n17811) );
  and2_0 U17278 ( .A(n17803), .B(n17804), .X(n17808) );
  o22ai_1 U17279 ( .A1(n17796), .A2(n17799), .B1(n17813), .B2(n17798), .Y(
        n17803) );
  o22ai_1 U17280 ( .A1(n11709), .A2(n11708), .B1(n11711), .B2(n17814), .Y(
        n17798) );
  and2_0 U17281 ( .A(n11708), .B(n11709), .X(n17814) );
  inv_1 U17282 ( .A(n17815), .Y(n11711) );
  o21ai_0 U17283 ( .A1(n12981), .A2(n17816), .B1(n12983), .Y(n17815) );
  nand2_1 U17284 ( .A(n17817), .B(n17818), .Y(n12983) );
  xor2_1 U17285 ( .A(n12726), .B(n12985), .X(n17816) );
  nor2_1 U17286 ( .A(n17818), .B(n17817), .Y(n12985) );
  xnor2_1 U17287 ( .A(n17819), .B(n10620), .Y(n17817) );
  xor2_1 U17288 ( .A(n17820), .B(n12959), .X(n17818) );
  o22ai_1 U17289 ( .A1(n16307), .A2(n17821), .B1(n17822), .B2(n17823), .Y(
        n17820) );
  inv_1 U17290 ( .A(n23763), .Y(n17823) );
  nor2_1 U17291 ( .A(n17824), .B(n11631), .Y(n17822) );
  and2_0 U17292 ( .A(n12994), .B(n17825), .X(n12981) );
  o22ai_1 U17293 ( .A1(n12993), .A2(n12992), .B1(n11079), .B2(n17826), .Y(
        n17825) );
  inv_1 U17294 ( .A(n11080), .Y(n17826) );
  nand2_1 U17295 ( .A(n17827), .B(n17828), .Y(n11080) );
  inv_1 U17296 ( .A(n12991), .Y(n11079) );
  nand2_1 U17297 ( .A(n11083), .B(n11082), .Y(n12991) );
  xor2_1 U17298 ( .A(n17829), .B(n17830), .X(n11082) );
  or2_0 U17299 ( .A(n17828), .B(n17827), .X(n17829) );
  mux2_1 U17300 ( .A0(n17831), .A1(n17832), .S(n17833), .X(n17827) );
  o21ai_0 U17301 ( .A1(n16870), .A2(n17834), .B1(n17835), .Y(n17832) );
  xor2_1 U17302 ( .A(n16870), .B(n17834), .X(n17831) );
  o22ai_1 U17303 ( .A1(n17003), .A2(n17836), .B1(n20744), .B2(n17837), .Y(
        n17828) );
  xor2_1 U17304 ( .A(n11413), .B(n17838), .X(n17837) );
  a21oi_1 U17305 ( .A1(n17839), .A2(n17069), .B1(n17840), .Y(n11083) );
  a21oi_1 U17306 ( .A1(n17841), .A2(n17068), .B1(n17067), .Y(n17840) );
  o21ai_0 U17307 ( .A1(n17003), .A2(n17842), .B1(n17843), .Y(n17067) );
  mux2i_1 U17308 ( .A0(n17844), .A1(n17838), .S(n17845), .Y(n17843) );
  and2_0 U17309 ( .A(n17003), .B(n17836), .X(n17838) );
  nor2_1 U17310 ( .A(n16277), .B(n17836), .Y(n17844) );
  xnor2_1 U17311 ( .A(n17845), .B(n17836), .Y(n17842) );
  xor2_1 U17312 ( .A(n17846), .B(outData[30]), .X(n17836) );
  xor2_1 U17313 ( .A(n20744), .B(n17340), .X(n17845) );
  inv_1 U17314 ( .A(n17841), .Y(n17069) );
  o21ai_0 U17315 ( .A1(n17847), .A2(n17080), .B1(n17081), .Y(n17841) );
  xnor2_1 U17316 ( .A(n11601), .B(n17848), .Y(n17081) );
  nor2_1 U17317 ( .A(n17849), .B(n17850), .Y(n17848) );
  o22ai_1 U17318 ( .A1(n17086), .A2(n17088), .B1(n17851), .B2(n17087), .Y(
        n17080) );
  xnor2_1 U17319 ( .A(n17852), .B(n17853), .Y(n17087) );
  xor2_1 U17320 ( .A(n12890), .B(n12485), .X(n17852) );
  and2_0 U17321 ( .A(n17086), .B(n17088), .X(n17851) );
  o22ai_1 U17322 ( .A1(n12901), .A2(n17854), .B1(n17855), .B2(n17856), .Y(
        n17088) );
  inv_1 U17323 ( .A(n23759), .Y(n17856) );
  nor2_1 U17324 ( .A(n17857), .B(n16637), .Y(n17855) );
  o22ai_1 U17325 ( .A1(n17858), .A2(n17859), .B1(n17057), .B2(n17061), .Y(
        n17086) );
  xor2_1 U17326 ( .A(n17860), .B(n17861), .X(n17061) );
  nor2_1 U17327 ( .A(n17059), .B(n17060), .Y(n17861) );
  inv_1 U17328 ( .A(n17859), .Y(n17059) );
  inv_1 U17329 ( .A(n17862), .Y(n17057) );
  o21ai_0 U17330 ( .A1(n17101), .A2(n17097), .B1(n17100), .Y(n17862) );
  nand2_1 U17331 ( .A(n17863), .B(n17864), .Y(n17100) );
  o22ai_1 U17332 ( .A1(n17107), .A2(n17106), .B1(n17108), .B2(n17865), .Y(
        n17097) );
  and2_0 U17333 ( .A(n17107), .B(n17106), .X(n17865) );
  a22oi_1 U17334 ( .A1(n17866), .A2(n17867), .B1(n17868), .B2(n23758), .Y(
        n17108) );
  o21ai_0 U17335 ( .A1(n16516), .A2(n17869), .B1(n17866), .Y(n17868) );
  inv_1 U17336 ( .A(n17870), .Y(n17867) );
  inv_1 U17337 ( .A(n17871), .Y(n17106) );
  a22oi_1 U17338 ( .A1(n17872), .A2(n17873), .B1(n17115), .B2(n17112), .Y(
        n17871) );
  mux2i_1 U17339 ( .A0(n17874), .A1(n17875), .S(n17598), .Y(n17112) );
  nor2_1 U17340 ( .A(n17092), .B(n17093), .Y(n17875) );
  xor2_1 U17341 ( .A(n17876), .B(n17877), .X(n17092) );
  o22ai_1 U17342 ( .A1(n17878), .A2(n17879), .B1(n17880), .B2(n17876), .Y(
        n17874) );
  xnor2_1 U17343 ( .A(n17881), .B(n17882), .Y(n17876) );
  xor2_1 U17344 ( .A(n23753), .B(n12297), .X(n17882) );
  nand2_1 U17345 ( .A(n17883), .B(n17884), .Y(n17881) );
  nor2_1 U17346 ( .A(n17877), .B(n17093), .Y(n17880) );
  inv_1 U17347 ( .A(n17093), .Y(n17879) );
  mux2i_1 U17348 ( .A0(n17885), .A1(n17886), .S(n11292), .Y(n17093) );
  nand2_1 U17349 ( .A(n17182), .B(n17887), .Y(n17886) );
  xor2_1 U17350 ( .A(n17888), .B(n17889), .X(n17182) );
  o22ai_1 U17351 ( .A1(n17183), .A2(n17889), .B1(n17890), .B2(n17888), .Y(
        n17885) );
  xnor2_1 U17352 ( .A(n16912), .B(n17891), .Y(n17888) );
  xor2_1 U17353 ( .A(n17892), .B(n17893), .X(n17891) );
  and2_0 U17354 ( .A(n17889), .B(n17183), .X(n17890) );
  o22ai_1 U17355 ( .A1(n17894), .A2(n16948), .B1(n23), .B2(n17895), .Y(n17889)
         );
  and2_0 U17356 ( .A(n16948), .B(n17894), .X(n17895) );
  inv_1 U17357 ( .A(n16916), .Y(n16948) );
  inv_1 U17358 ( .A(n17887), .Y(n17183) );
  o22ai_1 U17359 ( .A1(n17160), .A2(n17161), .B1(n17162), .B2(n17896), .Y(
        n17887) );
  and2_0 U17360 ( .A(n17161), .B(n17160), .X(n17896) );
  inv_1 U17361 ( .A(n17897), .Y(n17162) );
  o22ai_1 U17362 ( .A1(n16921), .A2(n17898), .B1(n17899), .B2(n17900), .Y(
        n17897) );
  inv_1 U17363 ( .A(n23683), .Y(n17900) );
  nor2_1 U17364 ( .A(n16583), .B(n17901), .Y(n17899) );
  xor2_1 U17365 ( .A(n23995), .B(n17898), .X(n17901) );
  o22ai_1 U17366 ( .A1(n17166), .A2(n17168), .B1(n17902), .B2(n17167), .Y(
        n17161) );
  o22ai_1 U17367 ( .A1(n16507), .A2(n17903), .B1(n17904), .B2(n17905), .Y(
        n17167) );
  inv_1 U17368 ( .A(n23756), .Y(n17905) );
  and2_0 U17369 ( .A(n17903), .B(n16507), .X(n17904) );
  and2_0 U17370 ( .A(n17168), .B(n17166), .X(n17902) );
  o21ai_0 U17371 ( .A1(n17178), .A2(n17172), .B1(n17177), .Y(n17168) );
  nand2_1 U17372 ( .A(n17906), .B(n17907), .Y(n17177) );
  mux2i_1 U17373 ( .A0(n17908), .A1(n17909), .S(n12984), .Y(n17172) );
  o22ai_1 U17374 ( .A1(n17910), .A2(n17911), .B1(n17912), .B2(n12659), .Y(
        n17909) );
  and2_0 U17375 ( .A(n17911), .B(n17910), .X(n17912) );
  nand2_1 U17376 ( .A(n12658), .B(n17913), .Y(n17908) );
  inv_1 U17377 ( .A(n12659), .Y(n17913) );
  xor2_1 U17378 ( .A(n17914), .B(n17915), .X(n12659) );
  o22ai_1 U17379 ( .A1(n16653), .A2(n16654), .B1(n16655), .B2(n17916), .Y(
        n17914) );
  and2_0 U17380 ( .A(n16654), .B(n16653), .X(n17916) );
  a22oi_1 U17381 ( .A1(n12650), .A2(n12648), .B1(n12647), .B2(n17917), .Y(
        n16655) );
  or2_0 U17382 ( .A(n12648), .B(n12650), .X(n17917) );
  nand2_1 U17383 ( .A(n17918), .B(n11584), .Y(n12647) );
  xor2_1 U17384 ( .A(n17919), .B(n11489), .X(n11584) );
  nand2_1 U17385 ( .A(n11585), .B(n11586), .Y(n17919) );
  inv_1 U17386 ( .A(n17920), .Y(n11586) );
  inv_1 U17387 ( .A(n17921), .Y(n11585) );
  xor2_1 U17388 ( .A(n12297), .B(n11583), .X(n17918) );
  a21oi_1 U17389 ( .A1(n17920), .A2(n17921), .B1(n11582), .Y(n11583) );
  o22ai_1 U17390 ( .A1(n17922), .A2(n16465), .B1(n17923), .B2(n16467), .Y(
        n11582) );
  xor2_1 U17391 ( .A(n17783), .B(n17924), .X(n16467) );
  xor2_1 U17392 ( .A(n2047), .B(n17925), .X(n17924) );
  and2_0 U17393 ( .A(n16465), .B(n17922), .X(n17923) );
  o22ai_1 U17394 ( .A1(n11136), .A2(n17926), .B1(n17927), .B2(n17928), .Y(
        n16465) );
  inv_1 U17395 ( .A(n23843), .Y(n17928) );
  and2_0 U17396 ( .A(n17926), .B(n11136), .X(n17927) );
  inv_1 U17397 ( .A(n16466), .Y(n17922) );
  o22ai_1 U17398 ( .A1(n16669), .A2(n16668), .B1(n17929), .B2(n17930), .Y(
        n16466) );
  and2_0 U17399 ( .A(n16668), .B(n16669), .X(n17930) );
  inv_1 U17400 ( .A(n16667), .Y(n17929) );
  o22ai_1 U17401 ( .A1(n16940), .A2(n17931), .B1(n21), .B2(n17932), .Y(n16667)
         );
  nor2_1 U17402 ( .A(n17933), .B(n12443), .Y(n17932) );
  inv_1 U17403 ( .A(n16940), .Y(n12443) );
  o22ai_1 U17404 ( .A1(n17934), .A2(n17935), .B1(n11042), .B2(n11039), .Y(
        n16668) );
  xnor2_1 U17405 ( .A(n17463), .B(n17936), .Y(n11039) );
  o21ai_0 U17406 ( .A1(n12454), .A2(n12455), .B1(n17937), .Y(n17936) );
  o21ai_0 U17407 ( .A1(n17938), .A2(n17939), .B1(n12449), .Y(n17937) );
  mux2i_1 U17408 ( .A0(n17940), .A1(n17941), .S(n32), .Y(n12449) );
  a21oi_1 U17409 ( .A1(n16674), .A2(n17942), .B1(n17943), .Y(n17941) );
  xor2_1 U17410 ( .A(n12731), .B(n17942), .X(n17940) );
  inv_1 U17411 ( .A(n12454), .Y(n17938) );
  inv_1 U17412 ( .A(n17939), .Y(n12455) );
  nor2_1 U17413 ( .A(n17944), .B(n11052), .Y(n17939) );
  xor2_1 U17414 ( .A(n16763), .B(n17945), .X(n11052) );
  nor2_1 U17415 ( .A(n17946), .B(n17947), .Y(n17945) );
  xor2_1 U17416 ( .A(n11168), .B(n17948), .X(n17944) );
  nor2_1 U17417 ( .A(n11051), .B(n11049), .Y(n17948) );
  xnor2_1 U17418 ( .A(n17949), .B(n12297), .Y(n11049) );
  o22ai_1 U17419 ( .A1(n16421), .A2(n16419), .B1(n17950), .B2(n16420), .Y(
        n17949) );
  xnor2_1 U17420 ( .A(n17951), .B(n17952), .Y(n16420) );
  o22ai_1 U17421 ( .A1(n16947), .A2(n17953), .B1(n23840), .B2(n17954), .Y(
        n17951) );
  xor2_1 U17422 ( .A(n17955), .B(n17956), .X(n17954) );
  nand2_1 U17423 ( .A(n16947), .B(n17953), .Y(n17956) );
  and2_0 U17424 ( .A(n16419), .B(n16421), .X(n17950) );
  o21ai_0 U17425 ( .A1(n11062), .A2(n11063), .B1(n17957), .Y(n16419) );
  xor2_1 U17426 ( .A(n11601), .B(n11061), .X(n17957) );
  o21ai_0 U17427 ( .A1(n11058), .A2(n11057), .B1(n11065), .Y(n11061) );
  xor2_1 U17428 ( .A(n17958), .B(n17959), .X(n11065) );
  nor2_1 U17429 ( .A(n17960), .B(n17961), .Y(n17959) );
  inv_1 U17430 ( .A(n11062), .Y(n17961) );
  xor2_1 U17431 ( .A(n17962), .B(n16750), .X(n11057) );
  nand3_1 U17432 ( .A(n17963), .B(n11063), .C(n11531), .Y(n17962) );
  inv_1 U17433 ( .A(n16686), .Y(n11058) );
  nand2_1 U17434 ( .A(n16687), .B(n17964), .Y(n16686) );
  xor2_1 U17435 ( .A(n23903), .B(n16690), .X(n17964) );
  a21oi_1 U17436 ( .A1(n11063), .A2(n17963), .B1(n11531), .Y(n16690) );
  nand2_1 U17437 ( .A(n16397), .B(n17965), .Y(n17963) );
  nor2_1 U17438 ( .A(n17966), .B(n17967), .Y(n16687) );
  inv_1 U17439 ( .A(n17960), .Y(n11063) );
  nor2_1 U17440 ( .A(n16397), .B(n17965), .Y(n17960) );
  o21ai_0 U17441 ( .A1(n16843), .A2(n17968), .B1(n17969), .Y(n17965) );
  xor2_1 U17442 ( .A(n17970), .B(n17971), .X(n17969) );
  nand2_1 U17443 ( .A(n17968), .B(n16843), .Y(n17971) );
  inv_1 U17444 ( .A(n42), .Y(n16397) );
  xor2_1 U17445 ( .A(n17972), .B(n17973), .X(n11062) );
  xor2_1 U17446 ( .A(n17953), .B(n16947), .X(n17973) );
  nand2_1 U17447 ( .A(n17974), .B(n17975), .Y(n17953) );
  o21ai_0 U17448 ( .A1(outData[7]), .A2(n17968), .B1(outData[8]), .Y(n17975)
         );
  xor2_1 U17449 ( .A(n17976), .B(n23840), .X(n17972) );
  xnor2_1 U17450 ( .A(n17793), .B(n17977), .Y(n16421) );
  xor2_1 U17451 ( .A(n2045), .B(n17978), .X(n17977) );
  and2_0 U17452 ( .A(n17946), .B(n17947), .X(n11051) );
  xor2_1 U17453 ( .A(n17979), .B(n17475), .X(n17947) );
  o22ai_1 U17454 ( .A1(n11120), .A2(n17980), .B1(n2045), .B2(n17981), .Y(
        n17979) );
  nor2_1 U17455 ( .A(n17978), .B(n17793), .Y(n17981) );
  inv_1 U17456 ( .A(n17978), .Y(n17980) );
  a21oi_1 U17457 ( .A1(n17974), .A2(outData[9]), .B1(n17982), .Y(n17978) );
  or3_1 U17458 ( .A(outData[8]), .B(outData[7]), .C(n17968), .X(n17974) );
  xor2_1 U17459 ( .A(n17983), .B(n17984), .X(n17946) );
  xor2_1 U17460 ( .A(n33), .B(n17985), .X(n17984) );
  xor2_1 U17461 ( .A(n16415), .B(n16902), .X(n17983) );
  o22ai_1 U17462 ( .A1(n16415), .A2(n17986), .B1(n33), .B2(n17987), .Y(n12454)
         );
  xor2_1 U17463 ( .A(n17988), .B(n17989), .X(n17987) );
  nor2_1 U17464 ( .A(n17985), .B(n16414), .Y(n17989) );
  inv_1 U17465 ( .A(n17985), .Y(n17986) );
  a21oi_1 U17466 ( .A1(n17990), .A2(outData[10]), .B1(n17991), .Y(n17985) );
  inv_1 U17467 ( .A(n17992), .Y(n17463) );
  xor2_1 U17468 ( .A(n12968), .B(n17993), .X(n11042) );
  nor2_1 U17469 ( .A(n11040), .B(n11041), .Y(n17993) );
  inv_1 U17470 ( .A(n11040), .Y(n17935) );
  xor2_1 U17471 ( .A(n17994), .B(n17931), .X(n11040) );
  inv_1 U17472 ( .A(n17933), .Y(n17931) );
  xor2_1 U17473 ( .A(n10617), .B(n17995), .X(n17933) );
  xor2_1 U17474 ( .A(n16940), .B(n21), .X(n17994) );
  inv_1 U17475 ( .A(n11041), .Y(n17934) );
  o22ai_1 U17476 ( .A1(n17996), .A2(n17997), .B1(n32), .B2(n17998), .Y(n11041)
         );
  xor2_1 U17477 ( .A(n17830), .B(n17943), .X(n17998) );
  nor2_1 U17478 ( .A(n16674), .B(n17942), .Y(n17943) );
  inv_1 U17479 ( .A(n17997), .Y(n17942) );
  o21ai_0 U17480 ( .A1(n17991), .A2(n10611), .B1(n17995), .Y(n17997) );
  xnor2_1 U17481 ( .A(n17999), .B(n16938), .Y(n16669) );
  xor2_1 U17482 ( .A(n17926), .B(n23843), .X(n17999) );
  nand2_1 U17483 ( .A(n18000), .B(n18001), .Y(n17926) );
  xor2_1 U17484 ( .A(n17403), .B(n18002), .X(n18000) );
  a21oi_1 U17485 ( .A1(n17995), .A2(outData[13]), .B1(n11173), .Y(n18002) );
  nor2_1 U17486 ( .A(n10617), .B(n12413), .Y(n11173) );
  o22ai_1 U17487 ( .A1(n17925), .A2(n17783), .B1(n2047), .B2(n18003), .Y(
        n17921) );
  and2_0 U17488 ( .A(n17783), .B(n17925), .X(n18003) );
  a21oi_1 U17489 ( .A1(n18001), .A2(outData[14]), .B1(n18004), .Y(n17925) );
  or3_1 U17490 ( .A(outData[13]), .B(outData[12]), .C(n17995), .X(n18001) );
  o21ai_0 U17491 ( .A1(n11130), .A2(n18005), .B1(n18006), .Y(n17920) );
  mux2i_1 U17492 ( .A0(n18007), .A1(n18008), .S(n18009), .Y(n18006) );
  nor2_1 U17493 ( .A(n18010), .B(n16933), .Y(n18008) );
  xor2_1 U17494 ( .A(n18010), .B(n18009), .X(n18005) );
  xor2_1 U17495 ( .A(n23845), .B(n12806), .X(n18009) );
  xnor2_1 U17496 ( .A(n18011), .B(n18012), .Y(n12648) );
  xor2_1 U17497 ( .A(n18013), .B(n18014), .X(n18012) );
  xor2_1 U17498 ( .A(n12640), .B(n18015), .X(n18011) );
  inv_1 U17499 ( .A(n12715), .Y(n12640) );
  nand2_1 U17500 ( .A(n18016), .B(n18017), .Y(n12650) );
  o21ai_0 U17501 ( .A1(n11130), .A2(n18018), .B1(n18019), .Y(n18017) );
  inv_1 U17502 ( .A(n23845), .Y(n18019) );
  xor2_1 U17503 ( .A(n17455), .B(n18010), .X(n18018) );
  inv_1 U17504 ( .A(n18020), .Y(n18010) );
  inv_1 U17505 ( .A(n11710), .Y(n17455) );
  xor2_1 U17506 ( .A(n18007), .B(n18021), .X(n18016) );
  nor2_1 U17507 ( .A(n18020), .B(n16933), .Y(n18007) );
  o21ai_0 U17508 ( .A1(n18022), .A2(n17633), .B1(n18023), .Y(n18020) );
  mux2i_1 U17509 ( .A0(n18024), .A1(n18025), .S(n16850), .Y(n18023) );
  nor2_1 U17510 ( .A(outData[15]), .B(n18004), .Y(n18024) );
  xor2_1 U17511 ( .A(n18004), .B(n18026), .X(n18022) );
  o22ai_1 U17512 ( .A1(n18027), .A2(n18028), .B1(n18029), .B2(n12705), .Y(
        n16654) );
  nor2_1 U17513 ( .A(n18027), .B(n18030), .Y(n18029) );
  inv_1 U17514 ( .A(n18031), .Y(n18027) );
  nor2_1 U17515 ( .A(n18032), .B(n18033), .Y(n16653) );
  a21oi_1 U17516 ( .A1(n18014), .A2(n12715), .B1(n18013), .Y(n18033) );
  inv_1 U17517 ( .A(n25), .Y(n18013) );
  xor2_1 U17518 ( .A(n18034), .B(n18035), .X(n18032) );
  nor2_1 U17519 ( .A(n12715), .B(n18014), .Y(n18035) );
  o21ai_0 U17520 ( .A1(n18025), .A2(n12310), .B1(n18036), .Y(n18014) );
  xor2_1 U17521 ( .A(n17911), .B(n17910), .X(n12658) );
  xor2_1 U17522 ( .A(n16482), .B(n18037), .X(n17910) );
  xnor2_1 U17523 ( .A(n23754), .B(n18038), .Y(n18037) );
  xor2_1 U17524 ( .A(n18039), .B(n18040), .X(n17911) );
  nand2_1 U17525 ( .A(n18031), .B(n18028), .Y(n18039) );
  or2_0 U17526 ( .A(n16925), .B(n18030), .X(n18028) );
  a21oi_1 U17527 ( .A1(n18041), .A2(n18042), .B1(n26), .Y(n18030) );
  nand3_1 U17528 ( .A(n18042), .B(n18041), .C(n26), .Y(n18031) );
  nand2_1 U17529 ( .A(outData[17]), .B(n18036), .Y(n18042) );
  xor2_1 U17530 ( .A(n11520), .B(n18043), .X(n17178) );
  nor2_1 U17531 ( .A(n17906), .B(n17907), .Y(n18043) );
  o22ai_1 U17532 ( .A1(n11386), .A2(n18038), .B1(n23754), .B2(n18044), .Y(
        n17907) );
  and2_0 U17533 ( .A(n18038), .B(n11386), .X(n18044) );
  o21ai_0 U17534 ( .A1(n18045), .A2(n11225), .B1(n18046), .Y(n18038) );
  xor2_1 U17535 ( .A(n18047), .B(n16507), .X(n17906) );
  xor2_1 U17536 ( .A(n17903), .B(n23756), .X(n18047) );
  o21ai_0 U17537 ( .A1(outData[19]), .A2(n10936), .B1(n18048), .Y(n17903) );
  xor2_1 U17538 ( .A(n18046), .B(n18049), .X(n18048) );
  nor2_1 U17539 ( .A(n18050), .B(n17051), .Y(n18049) );
  nand2_1 U17540 ( .A(n18045), .B(n11225), .Y(n18046) );
  inv_1 U17541 ( .A(n18050), .Y(n10936) );
  xnor2_1 U17542 ( .A(n18051), .B(n17898), .Y(n17166) );
  xor2_1 U17543 ( .A(n18052), .B(n18053), .X(n17898) );
  a21oi_1 U17544 ( .A1(outData[20]), .A2(n18054), .B1(n18055), .Y(n18053) );
  nand2_1 U17545 ( .A(n18056), .B(n11225), .Y(n18054) );
  xor2_1 U17546 ( .A(n16583), .B(n23683), .X(n18051) );
  xor2_1 U17547 ( .A(n18057), .B(n17894), .X(n17160) );
  xor2_1 U17548 ( .A(n18055), .B(n18058), .X(n17894) );
  xor2_1 U17549 ( .A(n11468), .B(n16493), .X(n18058) );
  xor2_1 U17550 ( .A(n23), .B(n16916), .X(n18057) );
  inv_1 U17551 ( .A(n17877), .Y(n17878) );
  nor2_1 U17552 ( .A(n18059), .B(n18060), .Y(n17877) );
  a21oi_1 U17553 ( .A1(n17893), .A2(n16561), .B1(n17892), .Y(n18060) );
  inv_1 U17554 ( .A(n23757), .Y(n17892) );
  inv_1 U17555 ( .A(n16912), .Y(n16561) );
  xor2_1 U17556 ( .A(n18061), .B(n17611), .X(n18059) );
  nor2_1 U17557 ( .A(n18062), .B(n17893), .Y(n18061) );
  nand2_1 U17558 ( .A(n18063), .B(n18064), .Y(n17893) );
  o21ai_0 U17559 ( .A1(outData[21]), .A2(n18065), .B1(outData[22]), .Y(n18063)
         );
  inv_1 U17560 ( .A(n18055), .Y(n18065) );
  xor2_1 U17561 ( .A(n16912), .B(n18066), .X(n18062) );
  xnor2_1 U17562 ( .A(n18067), .B(n18068), .Y(n17115) );
  nand2_1 U17563 ( .A(n17113), .B(n17114), .Y(n18067) );
  inv_1 U17564 ( .A(n17872), .Y(n17113) );
  inv_1 U17565 ( .A(n17114), .Y(n17873) );
  xor2_1 U17566 ( .A(n16520), .B(n18069), .X(n17114) );
  nor2_1 U17567 ( .A(n18070), .B(n18071), .Y(n18069) );
  inv_1 U17568 ( .A(n18072), .Y(n18071) );
  o21ai_0 U17569 ( .A1(n23753), .A2(n18073), .B1(n18074), .Y(n17872) );
  xnor2_1 U17570 ( .A(n16931), .B(n17884), .Y(n18074) );
  nand2_1 U17571 ( .A(n18075), .B(n16550), .Y(n17884) );
  xor2_1 U17572 ( .A(n18076), .B(n11284), .X(n18075) );
  xor2_1 U17573 ( .A(n18077), .B(n17883), .X(n18073) );
  nand2_1 U17574 ( .A(n18078), .B(n17766), .Y(n17883) );
  xor2_1 U17575 ( .A(n11622), .B(n18076), .X(n18078) );
  nand2_1 U17576 ( .A(n18079), .B(n18080), .Y(n18076) );
  xor2_1 U17577 ( .A(n17133), .B(n18081), .X(n18079) );
  nand2_1 U17578 ( .A(outData[23]), .B(n18064), .Y(n18081) );
  o21ai_0 U17579 ( .A1(n18082), .A2(n16520), .B1(n18072), .Y(n17107) );
  o211ai_1 U17580 ( .A1(n18083), .A2(n17709), .B1(n16906), .C1(n18084), .Y(
        n18072) );
  inv_1 U17581 ( .A(n23682), .Y(n16520) );
  xor2_1 U17582 ( .A(n17644), .B(n18070), .X(n18082) );
  and2_0 U17583 ( .A(n16542), .B(n18085), .X(n18070) );
  o21ai_0 U17584 ( .A1(n18083), .A2(n17709), .B1(n18084), .Y(n18085) );
  xor2_1 U17585 ( .A(n18086), .B(n18087), .X(n17101) );
  nor2_1 U17586 ( .A(n17863), .B(n17864), .Y(n18087) );
  xor2_1 U17587 ( .A(n18088), .B(n17830), .X(n17864) );
  nand2_1 U17588 ( .A(n17870), .B(n17866), .Y(n18088) );
  nand2_1 U17589 ( .A(n17869), .B(n16516), .Y(n17866) );
  o21ai_0 U17590 ( .A1(n17869), .A2(n16516), .B1(n16629), .Y(n17870) );
  inv_1 U17591 ( .A(n23758), .Y(n16629) );
  a21oi_1 U17592 ( .A1(n18084), .A2(outData[25]), .B1(n18089), .Y(n17869) );
  xor2_1 U17593 ( .A(n16625), .B(n18090), .X(n17863) );
  xor2_1 U17594 ( .A(n24), .B(n18091), .X(n18090) );
  xor2_1 U17595 ( .A(n12901), .B(n18092), .X(n17859) );
  xor2_1 U17596 ( .A(n23759), .B(n17857), .X(n18092) );
  inv_1 U17597 ( .A(n17854), .Y(n17857) );
  o21ai_0 U17598 ( .A1(n12412), .A2(n18093), .B1(n18094), .Y(n17854) );
  mux2i_1 U17599 ( .A0(n18095), .A1(n18096), .S(n13351), .Y(n18094) );
  and2_0 U17600 ( .A(n18097), .B(n12412), .X(n18096) );
  xor2_1 U17601 ( .A(n13368), .B(n18097), .X(n18093) );
  inv_1 U17602 ( .A(n17060), .Y(n17858) );
  nand2_1 U17603 ( .A(n18098), .B(n18099), .Y(n17060) );
  o21ai_0 U17604 ( .A1(n18091), .A2(n16625), .B1(n24), .Y(n18099) );
  inv_1 U17605 ( .A(n18100), .Y(n18091) );
  xor2_1 U17606 ( .A(n16757), .B(n18101), .X(n18098) );
  nor2_1 U17607 ( .A(n12907), .B(n18100), .Y(n18101) );
  o21ai_0 U17608 ( .A1(n18089), .A2(n17711), .B1(n18097), .Y(n18100) );
  inv_1 U17609 ( .A(n17082), .Y(n17847) );
  nand2_1 U17610 ( .A(n17849), .B(n17850), .Y(n17082) );
  o22ai_1 U17611 ( .A1(n16894), .A2(n17853), .B1(n12485), .B2(n18102), .Y(
        n17850) );
  and2_0 U17612 ( .A(n16894), .B(n17853), .X(n18102) );
  xnor2_1 U17613 ( .A(n18103), .B(n18095), .Y(n17853) );
  xor2_1 U17614 ( .A(n11336), .B(outData[28]), .X(n18103) );
  xor2_1 U17615 ( .A(n18104), .B(n16280), .X(n17849) );
  o21ai_0 U17616 ( .A1(n16882), .A2(n18105), .B1(n18106), .Y(n18104) );
  inv_1 U17617 ( .A(n17068), .Y(n17839) );
  mux2i_1 U17618 ( .A0(n18107), .A1(n18108), .S(n23903), .Y(n17068) );
  a22oi_1 U17619 ( .A1(n18106), .A2(n16280), .B1(n18109), .B2(n18110), .Y(
        n18108) );
  inv_1 U17620 ( .A(n23760), .Y(n16280) );
  nand2_1 U17621 ( .A(n18105), .B(n16882), .Y(n18106) );
  nor2_1 U17622 ( .A(n18105), .B(n18111), .Y(n18107) );
  inv_1 U17623 ( .A(n18109), .Y(n18105) );
  xor2_1 U17624 ( .A(n18112), .B(n18015), .X(n18109) );
  o211ai_1 U17625 ( .A1(n18095), .A2(n11498), .B1(n11497), .C1(n18113), .Y(
        n18112) );
  nand2_1 U17626 ( .A(outData[29]), .B(outData[28]), .Y(n11497) );
  xnor2_1 U17627 ( .A(n11185), .B(n18114), .Y(n12994) );
  and2_0 U17628 ( .A(n12992), .B(n12993), .X(n18114) );
  xor2_1 U17629 ( .A(n11631), .B(n18115), .X(n12993) );
  xor2_1 U17630 ( .A(n23763), .B(n17824), .X(n18115) );
  nand2_1 U17631 ( .A(n18116), .B(n18117), .Y(n12992) );
  o21ai_0 U17632 ( .A1(n16870), .A2(n17834), .B1(n17833), .Y(n18117) );
  inv_1 U17633 ( .A(n23693), .Y(n17833) );
  xor2_1 U17634 ( .A(n17066), .B(n17835), .X(n18116) );
  nand2_1 U17635 ( .A(n17834), .B(n16870), .Y(n17835) );
  inv_1 U17636 ( .A(n16872), .Y(n16870) );
  xor2_1 U17637 ( .A(n18118), .B(n18119), .X(n17834) );
  a21oi_1 U17638 ( .A1(n18120), .A2(n17846), .B1(n17824), .Y(n18119) );
  inv_1 U17639 ( .A(n18113), .Y(n17846) );
  nand2_1 U17640 ( .A(n18121), .B(n18122), .Y(n11708) );
  o21ai_0 U17641 ( .A1(n17824), .A2(n11763), .B1(n10620), .Y(n18122) );
  mux2i_1 U17642 ( .A0(n17819), .A1(n18123), .S(n16773), .Y(n18121) );
  nor2_1 U17643 ( .A(n16314), .B(n17821), .Y(n18123) );
  xor2_1 U17644 ( .A(n11763), .B(n17824), .X(n17819) );
  inv_1 U17645 ( .A(n17821), .Y(n17824) );
  o21ai_0 U17646 ( .A1(outData[30]), .A2(n18113), .B1(n18124), .Y(n17821) );
  nand3_1 U17647 ( .A(n10612), .B(n11498), .C(n18095), .Y(n18113) );
  nor2_1 U17648 ( .A(n18097), .B(outData[27]), .Y(n18095) );
  nand2_1 U17649 ( .A(n18089), .B(n17711), .Y(n18097) );
  nor2_1 U17650 ( .A(n18084), .B(outData[25]), .Y(n18089) );
  xnor2_1 U17651 ( .A(n18125), .B(n18126), .Y(n18084) );
  nor2_1 U17652 ( .A(outData[24]), .B(n18080), .Y(n18126) );
  inv_1 U17653 ( .A(n18083), .Y(n18080) );
  xor2_1 U17654 ( .A(n18127), .B(n18128), .X(n18083) );
  or2_0 U17655 ( .A(n18064), .B(outData[23]), .X(n18127) );
  nand3_1 U17656 ( .A(n12426), .B(n11468), .C(n18055), .Y(n18064) );
  xor2_1 U17657 ( .A(n18129), .B(n18130), .X(n18055) );
  and2_0 U17658 ( .A(n18056), .B(n18131), .X(n18130) );
  nor2_1 U17659 ( .A(n18041), .B(outData[19]), .Y(n18056) );
  inv_1 U17660 ( .A(n18045), .Y(n18041) );
  nor2_1 U17661 ( .A(n18036), .B(outData[17]), .Y(n18045) );
  nand2_1 U17662 ( .A(n18025), .B(n12310), .Y(n18036) );
  and2_0 U17663 ( .A(n18004), .B(n17633), .X(n18025) );
  nor3_1 U17664 ( .A(n17995), .B(outData[13]), .C(n18132), .Y(n18004) );
  xnor2_1 U17665 ( .A(n18133), .B(n11570), .Y(n17995) );
  nand2_1 U17666 ( .A(n17991), .B(n10611), .Y(n18133) );
  nor2_1 U17667 ( .A(n17990), .B(outData[10]), .Y(n17991) );
  inv_1 U17668 ( .A(n17982), .Y(n17990) );
  nor3_1 U17669 ( .A(n17968), .B(outData[8]), .C(n18134), .Y(n17982) );
  xnor2_1 U17670 ( .A(n18135), .B(n18136), .Y(n17968) );
  nand4_1 U17671 ( .A(n18137), .B(n18138), .C(n12440), .D(n10604), .Y(n18135)
         );
  xor2_1 U17672 ( .A(n16763), .B(n18139), .X(n18137) );
  nor3_1 U17673 ( .A(outData[2]), .B(outData[6]), .C(outData[3]), .Y(n18139)
         );
  xnor2_1 U17674 ( .A(n18140), .B(n13031), .Y(n11709) );
  xor2_1 U17675 ( .A(n10620), .B(n12351), .X(n18140) );
  and2_0 U17676 ( .A(n17799), .B(n17796), .X(n17813) );
  xnor2_1 U17677 ( .A(n11755), .B(n18141), .Y(n17799) );
  xor2_1 U17678 ( .A(n23875), .B(n12351), .X(n18141) );
  xor2_1 U17679 ( .A(n17031), .B(n18142), .X(n17796) );
  a21oi_1 U17680 ( .A1(n16863), .A2(n17810), .B1(n18143), .Y(n18142) );
  a21oi_1 U17681 ( .A1(n12351), .A2(n13031), .B1(n10620), .Y(n18143) );
  inv_1 U17682 ( .A(n12351), .Y(n17810) );
  xor2_1 U17683 ( .A(n18144), .B(n16229), .X(n17804) );
  xor2_1 U17684 ( .A(n10811), .B(n23875), .X(n18144) );
  nand2_1 U17685 ( .A(n18145), .B(n10815), .Y(n17806) );
  nand2_1 U17686 ( .A(n18146), .B(n18147), .Y(n10815) );
  inv_1 U17687 ( .A(n10816), .Y(n18145) );
  xor2_1 U17688 ( .A(n16464), .B(n18148), .X(n10816) );
  nor2_1 U17689 ( .A(n18146), .B(n18147), .Y(n18148) );
  o22ai_1 U17690 ( .A1(n16226), .A2(n10811), .B1(n23875), .B2(n18149), .Y(
        n18147) );
  nor2_1 U17691 ( .A(n23765), .B(n16229), .Y(n18149) );
  inv_1 U17692 ( .A(n23765), .Y(n10811) );
  xor2_1 U17693 ( .A(n10810), .B(n18150), .X(n18146) );
  xor2_1 U17694 ( .A(n20745), .B(n23765), .X(n18150) );
  nand2_1 U17695 ( .A(n18151), .B(n11593), .Y(n10147) );
  inv_1 U17696 ( .A(n10802), .Y(n11593) );
  nand2_1 U17697 ( .A(n18152), .B(n15868), .Y(n10802) );
  inv_1 U17698 ( .A(n15853), .Y(n15868) );
  nor2_1 U17699 ( .A(n11703), .B(n24062), .Y(n15853) );
  mux2i_1 U17700 ( .A0(n18153), .A1(n18154), .S(n10819), .Y(n18151) );
  nand2_1 U17701 ( .A(inData[2]), .B(n18155), .Y(n18154) );
  xor2_1 U17702 ( .A(n66), .B(n10823), .X(n18155) );
  nor2_1 U17703 ( .A(n11508), .B(n23721), .Y(n10823) );
  inv_1 U17704 ( .A(n23769), .Y(n11508) );
  xor2_1 U17705 ( .A(n18156), .B(n10827), .X(n18153) );
  inv_1 U17706 ( .A(n10848), .Y(n10827) );
  xor2_1 U17707 ( .A(n18157), .B(n18158), .X(n10848) );
  xor2_1 U17708 ( .A(n12380), .B(n18159), .X(n18158) );
  a21oi_1 U17709 ( .A1(n18160), .A2(n18161), .B1(n18162), .Y(n18159) );
  inv_1 U17710 ( .A(n18163), .Y(n18161) );
  xor2_1 U17711 ( .A(n17338), .B(n18164), .X(n18160) );
  a21oi_1 U17712 ( .A1(n18165), .A2(n18166), .B1(n10826), .Y(n18164) );
  xor2_1 U17713 ( .A(n10828), .B(n23680), .X(n18156) );
  o22ai_1 U17714 ( .A1(n18167), .A2(n11528), .B1(n18168), .B2(n18169), .Y(
        n10828) );
  inv_1 U17715 ( .A(n23770), .Y(n18169) );
  and2_0 U17716 ( .A(n11528), .B(n18167), .X(n18168) );
  o22ai_1 U17717 ( .A1(n23721), .A2(n10821), .B1(n10819), .B2(n18170), .Y(
        n10146) );
  xor2_1 U17718 ( .A(n11528), .B(n18171), .X(n18170) );
  xor2_1 U17719 ( .A(n23770), .B(n18167), .X(n18171) );
  a22oi_1 U17720 ( .A1(n11715), .A2(n11716), .B1(n18172), .B2(n15), .Y(n18167)
         );
  or2_0 U17721 ( .A(n11716), .B(n11715), .X(n18172) );
  a21oi_1 U17722 ( .A1(n11602), .A2(n11603), .B1(n18173), .Y(n11716) );
  inv_1 U17723 ( .A(n18174), .Y(n18173) );
  o21ai_0 U17724 ( .A1(n11603), .A2(n11602), .B1(n23772), .Y(n18174) );
  xnor2_1 U17725 ( .A(n18175), .B(n18176), .Y(n11603) );
  xor2_1 U17726 ( .A(n18177), .B(n18178), .X(n18176) );
  nand2_1 U17727 ( .A(n18179), .B(n18180), .Y(n18177) );
  o32ai_1 U17728 ( .A1(n18181), .A2(n18182), .A3(n18183), .B1(n18183), .B2(
        n10826), .Y(n18180) );
  xor2_1 U17729 ( .A(n18184), .B(n12380), .X(n18175) );
  o22ai_1 U17730 ( .A1(n11727), .A2(n17124), .B1(n16), .B2(n18185), .Y(n11602)
         );
  and2_0 U17731 ( .A(n17124), .B(n11727), .X(n18185) );
  o22ai_1 U17732 ( .A1(n12999), .A2(n12998), .B1(n18186), .B2(n18187), .Y(
        n17124) );
  inv_1 U17733 ( .A(n23681), .Y(n18187) );
  nor2_1 U17734 ( .A(n13006), .B(n18188), .Y(n18186) );
  inv_1 U17735 ( .A(n12998), .Y(n13006) );
  xor2_1 U17736 ( .A(n18189), .B(n18190), .X(n12998) );
  xor2_1 U17737 ( .A(n18191), .B(n18192), .X(n18190) );
  a21oi_1 U17738 ( .A1(n18193), .A2(n10826), .B1(n18182), .Y(n18191) );
  xor2_1 U17739 ( .A(n11520), .B(n12380), .X(n18189) );
  inv_1 U17740 ( .A(n18188), .Y(n12999) );
  o22ai_1 U17741 ( .A1(n11089), .A2(n11092), .B1(n18194), .B2(n11091), .Y(
        n18188) );
  inv_1 U17742 ( .A(n23773), .Y(n11091) );
  and2_0 U17743 ( .A(n11092), .B(n11089), .X(n18194) );
  o22ai_1 U17744 ( .A1(n17138), .A2(n17139), .B1(n18195), .B2(n17075), .Y(
        n11092) );
  inv_1 U17745 ( .A(n23774), .Y(n17075) );
  and2_0 U17746 ( .A(n17139), .B(n17138), .X(n18195) );
  o22ai_1 U17747 ( .A1(n17146), .A2(n17145), .B1(n23775), .B2(n18196), .Y(
        n17139) );
  and2_0 U17748 ( .A(n17145), .B(n17146), .X(n18196) );
  o21ai_0 U17749 ( .A1(n17150), .A2(n10632), .B1(n18197), .Y(n17145) );
  xor2_1 U17750 ( .A(n14685), .B(n18198), .X(n18197) );
  nand2_1 U17751 ( .A(n17148), .B(n17153), .Y(n18198) );
  nand2_1 U17752 ( .A(n17150), .B(n10632), .Y(n17153) );
  o22ai_1 U17753 ( .A1(n17132), .A2(n18199), .B1(n18200), .B2(n17070), .Y(
        n17148) );
  inv_1 U17754 ( .A(n17), .Y(n17070) );
  nor2_1 U17755 ( .A(n17131), .B(n17689), .Y(n18200) );
  inv_1 U17756 ( .A(n17131), .Y(n18199) );
  a22oi_1 U17757 ( .A1(n17682), .A2(n17194), .B1(n18201), .B2(n23778), .Y(
        n17131) );
  or2_0 U17758 ( .A(n17194), .B(n17682), .X(n18201) );
  mux2i_1 U17759 ( .A0(n18202), .A1(n18203), .S(n18204), .Y(n17194) );
  o22ai_1 U17760 ( .A1(n16982), .A2(n18205), .B1(n18206), .B2(n10643), .Y(
        n18203) );
  nor2_1 U17761 ( .A(n17670), .B(n18207), .Y(n18206) );
  inv_1 U17762 ( .A(n17670), .Y(n18205) );
  inv_1 U17763 ( .A(n18207), .Y(n16982) );
  nand2_1 U17764 ( .A(n16981), .B(n18207), .Y(n18202) );
  o22ai_1 U17765 ( .A1(n16975), .A2(n16977), .B1(n18208), .B2(n10634), .Y(
        n18207) );
  and2_0 U17766 ( .A(n16977), .B(n16975), .X(n18208) );
  o221ai_1 U17767 ( .A1(n17036), .A2(n17187), .B1(n18209), .B2(n17189), .C1(
        n18210), .Y(n16977) );
  o21ai_0 U17768 ( .A1(n18211), .A2(n18212), .B1(n23783), .Y(n18210) );
  inv_1 U17769 ( .A(n17189), .Y(n18212) );
  nor2_1 U17770 ( .A(n18213), .B(n18209), .Y(n18211) );
  o22ai_1 U17771 ( .A1(n17198), .A2(n17200), .B1(n18214), .B2(n17157), .Y(
        n17189) );
  inv_1 U17772 ( .A(n23780), .Y(n17157) );
  and2_0 U17773 ( .A(n17200), .B(n17198), .X(n18214) );
  o22ai_1 U17774 ( .A1(n17205), .A2(n17638), .B1(n18215), .B2(n18216), .Y(
        n17200) );
  inv_1 U17775 ( .A(n23781), .Y(n18216) );
  and2_0 U17776 ( .A(n17205), .B(n17638), .X(n18215) );
  o21ai_0 U17777 ( .A1(n12302), .A2(n18217), .B1(n18218), .Y(n17638) );
  mux2i_1 U17778 ( .A0(n18219), .A1(n18220), .S(n18221), .Y(n18218) );
  nor2_1 U17779 ( .A(n18222), .B(n15931), .Y(n18220) );
  xor2_1 U17780 ( .A(n18223), .B(n18224), .X(n18217) );
  o21ai_0 U17781 ( .A1(n23696), .A2(n17216), .B1(n18225), .Y(n17205) );
  xor2_1 U17782 ( .A(n12939), .B(n18226), .X(n18225) );
  nand2_1 U17783 ( .A(n17215), .B(n17217), .Y(n18226) );
  nand2_1 U17784 ( .A(n23696), .B(n17216), .Y(n17217) );
  xor2_1 U17785 ( .A(n18227), .B(n12297), .X(n17215) );
  o22ai_1 U17786 ( .A1(n17222), .A2(n17220), .B1(n23691), .B2(n18228), .Y(
        n18227) );
  and2_0 U17787 ( .A(n17220), .B(n17222), .X(n18228) );
  xor2_1 U17788 ( .A(n18229), .B(n23959), .X(n17220) );
  nand2_1 U17789 ( .A(n18230), .B(n18231), .Y(n18229) );
  inv_1 U17790 ( .A(n18232), .Y(n17222) );
  o22ai_1 U17791 ( .A1(n12665), .A2(n18233), .B1(n18234), .B2(n12666), .Y(
        n18232) );
  inv_1 U17792 ( .A(n23782), .Y(n12666) );
  nor2_1 U17793 ( .A(n12667), .B(n17493), .Y(n18234) );
  inv_1 U17794 ( .A(n18233), .Y(n12667) );
  o22ai_1 U17795 ( .A1(n12671), .A2(n12673), .B1(n12430), .B2(n18235), .Y(
        n18233) );
  and2_0 U17796 ( .A(n12673), .B(n12671), .X(n18235) );
  o22ai_1 U17797 ( .A1(n18236), .A2(n17503), .B1(n18237), .B2(n16706), .Y(
        n12673) );
  inv_1 U17798 ( .A(n18), .Y(n16706) );
  nor2_1 U17799 ( .A(n16705), .B(n16704), .Y(n18237) );
  inv_1 U17800 ( .A(n16705), .Y(n17503) );
  xor2_1 U17801 ( .A(n18238), .B(n18239), .X(n16705) );
  xor2_1 U17802 ( .A(n18240), .B(n18241), .X(n18239) );
  xor2_1 U17803 ( .A(n18026), .B(n1965), .X(n18238) );
  inv_1 U17804 ( .A(n16704), .Y(n18236) );
  o22ai_1 U17805 ( .A1(n17618), .A2(n11591), .B1(n18242), .B2(n18243), .Y(
        n16704) );
  inv_1 U17806 ( .A(n55), .Y(n18243) );
  and2_0 U17807 ( .A(n11591), .B(n17618), .X(n18242) );
  o22ai_1 U17808 ( .A1(n17529), .A2(n12678), .B1(n18244), .B2(n12447), .Y(
        n11591) );
  inv_1 U17809 ( .A(n23711), .Y(n12447) );
  and2_0 U17810 ( .A(n12678), .B(n17529), .X(n18244) );
  o22ai_1 U17811 ( .A1(n18245), .A2(n18246), .B1(n18247), .B2(n12656), .Y(
        n12678) );
  inv_1 U17812 ( .A(n23848), .Y(n12656) );
  nor2_1 U17813 ( .A(n16719), .B(n16721), .Y(n18247) );
  inv_1 U17814 ( .A(n16719), .Y(n18246) );
  xor2_1 U17815 ( .A(n18248), .B(n23981), .X(n16719) );
  nand2_1 U17816 ( .A(n18249), .B(n18250), .Y(n18248) );
  xor2_1 U17817 ( .A(n18125), .B(n18251), .X(n18249) );
  inv_1 U17818 ( .A(n16721), .Y(n18245) );
  o22ai_1 U17819 ( .A1(n16710), .A2(n16711), .B1(n18252), .B2(n11046), .Y(
        n16721) );
  inv_1 U17820 ( .A(n12517), .Y(n11046) );
  and2_0 U17821 ( .A(n16711), .B(n16710), .X(n18252) );
  o22ai_1 U17822 ( .A1(n18253), .A2(n17548), .B1(n18254), .B2(n12465), .Y(
        n16711) );
  inv_1 U17823 ( .A(n23850), .Y(n12465) );
  nor2_1 U17824 ( .A(n16698), .B(n16699), .Y(n18254) );
  inv_1 U17825 ( .A(n17548), .Y(n16698) );
  xnor2_1 U17826 ( .A(n18255), .B(n18256), .Y(n17548) );
  xor2_1 U17827 ( .A(n16453), .B(n18257), .X(n18255) );
  inv_1 U17828 ( .A(n16699), .Y(n18253) );
  o22ai_1 U17829 ( .A1(n16714), .A2(n17603), .B1(n18258), .B2(n16685), .Y(
        n16699) );
  inv_1 U17830 ( .A(n23878), .Y(n16685) );
  nor2_1 U17831 ( .A(n16716), .B(n18259), .Y(n18258) );
  inv_1 U17832 ( .A(n16714), .Y(n18259) );
  inv_1 U17833 ( .A(n16716), .Y(n17603) );
  xor2_1 U17834 ( .A(n18260), .B(n18261), .X(n16716) );
  xor2_1 U17835 ( .A(n18262), .B(n17525), .X(n18261) );
  nand2_1 U17836 ( .A(n18263), .B(n18264), .Y(n18260) );
  inv_1 U17837 ( .A(n18265), .Y(n18263) );
  xor2_1 U17838 ( .A(n18266), .B(n16850), .X(n16714) );
  o22ai_1 U17839 ( .A1(n18267), .A2(n17587), .B1(n2046), .B2(n18268), .Y(
        n18266) );
  nor2_1 U17840 ( .A(n16695), .B(n16694), .Y(n18268) );
  inv_1 U17841 ( .A(n16695), .Y(n17587) );
  xor2_1 U17842 ( .A(n18269), .B(n12388), .X(n16695) );
  nand2_1 U17843 ( .A(n18270), .B(n18271), .Y(n18269) );
  inv_1 U17844 ( .A(n16694), .Y(n18267) );
  o21ai_0 U17845 ( .A1(n23877), .A2(n11070), .B1(n18272), .Y(n16694) );
  xor2_1 U17846 ( .A(n17338), .B(n18273), .X(n18272) );
  a21oi_1 U17847 ( .A1(n23877), .A2(n11070), .B1(n11071), .Y(n18273) );
  inv_1 U17848 ( .A(n16724), .Y(n11071) );
  nor2_1 U17849 ( .A(n16723), .B(n20), .Y(n16724) );
  xor2_1 U17850 ( .A(n18274), .B(n18275), .X(n16723) );
  nand2_1 U17851 ( .A(n18276), .B(n18277), .Y(n18274) );
  inv_1 U17852 ( .A(n16627), .Y(n17338) );
  inv_1 U17853 ( .A(n17565), .Y(n11070) );
  xor2_1 U17854 ( .A(n15972), .B(n18278), .X(n17565) );
  a21oi_1 U17855 ( .A1(n18279), .A2(n16818), .B1(n18280), .Y(n18278) );
  xor2_1 U17856 ( .A(n17774), .B(n18281), .X(n18280) );
  inv_1 U17857 ( .A(n17541), .Y(n16710) );
  xnor2_1 U17858 ( .A(n18282), .B(n18283), .Y(n17541) );
  xor2_1 U17859 ( .A(n18284), .B(n12394), .X(n18282) );
  inv_1 U17860 ( .A(n12676), .Y(n17529) );
  xor2_1 U17861 ( .A(n18285), .B(n12392), .X(n12676) );
  nand2_1 U17862 ( .A(n18286), .B(n18287), .Y(n18285) );
  xor2_1 U17863 ( .A(n18288), .B(n18289), .X(n17618) );
  xor2_1 U17864 ( .A(n18290), .B(n18291), .X(n18289) );
  inv_1 U17865 ( .A(n18292), .Y(n18291) );
  xor2_1 U17866 ( .A(n16510), .B(n12297), .X(n18288) );
  xor2_1 U17867 ( .A(n18293), .B(n18294), .X(n12671) );
  xor2_1 U17868 ( .A(n15902), .B(n18295), .X(n18294) );
  inv_1 U17869 ( .A(n17493), .Y(n12665) );
  xor2_1 U17870 ( .A(n18296), .B(n18297), .X(n17493) );
  xor2_1 U17871 ( .A(n23958), .B(n18298), .X(n18297) );
  xor2_1 U17872 ( .A(n18299), .B(n16524), .X(n17216) );
  nand2_1 U17873 ( .A(n18300), .B(n18301), .Y(n18299) );
  inv_1 U17874 ( .A(n18302), .Y(n18301) );
  xnor2_1 U17875 ( .A(n18303), .B(n18304), .Y(n17198) );
  xor2_1 U17876 ( .A(n18305), .B(n18306), .X(n18304) );
  xor2_1 U17877 ( .A(n18209), .B(n23783), .X(n17187) );
  inv_1 U17878 ( .A(n17467), .Y(n18209) );
  xnor2_1 U17879 ( .A(n18307), .B(n18308), .Y(n17467) );
  xor2_1 U17880 ( .A(n18309), .B(n16611), .X(n18307) );
  xor2_1 U17881 ( .A(n18310), .B(n18311), .X(n16975) );
  xor2_1 U17882 ( .A(n18312), .B(n12299), .X(n18310) );
  xor2_1 U17883 ( .A(n17670), .B(n23784), .X(n16981) );
  xor2_1 U17884 ( .A(n18313), .B(n18314), .X(n17670) );
  xor2_1 U17885 ( .A(n18315), .B(n11048), .X(n18314) );
  xor2_1 U17886 ( .A(n18316), .B(n23951), .X(n18313) );
  inv_1 U17887 ( .A(n17195), .Y(n17682) );
  xor2_1 U17888 ( .A(n18317), .B(n18318), .X(n17195) );
  xor2_1 U17889 ( .A(n23903), .B(n12320), .X(n18318) );
  xor2_1 U17890 ( .A(n18319), .B(n18320), .X(n18317) );
  inv_1 U17891 ( .A(n17689), .Y(n17132) );
  o22ai_1 U17892 ( .A1(n18321), .A2(n18322), .B1(n23938), .B2(n18323), .Y(
        n17689) );
  and2_0 U17893 ( .A(n18324), .B(n18325), .X(n18323) );
  inv_1 U17894 ( .A(n18324), .Y(n18321) );
  inv_1 U17895 ( .A(n17453), .Y(n17150) );
  xor2_1 U17896 ( .A(n18326), .B(n18327), .X(n17453) );
  xor2_1 U17897 ( .A(n10607), .B(n11574), .X(n18327) );
  xor2_1 U17898 ( .A(n18328), .B(n18329), .X(n18326) );
  xor2_1 U17899 ( .A(n18330), .B(n23949), .X(n17146) );
  nand2_1 U17900 ( .A(n18331), .B(n18332), .Y(n18330) );
  xnor2_1 U17901 ( .A(n18333), .B(n18334), .Y(n17138) );
  xor2_1 U17902 ( .A(n18335), .B(n18336), .X(n18334) );
  xor2_1 U17903 ( .A(n10826), .B(n18068), .X(n18333) );
  xor2_1 U17904 ( .A(n18337), .B(n18338), .X(n11089) );
  xor2_1 U17905 ( .A(n10826), .B(n16742), .X(n18338) );
  xor2_1 U17906 ( .A(n18193), .B(n18339), .X(n18337) );
  xor2_1 U17907 ( .A(n18340), .B(n18341), .X(n11727) );
  xor2_1 U17908 ( .A(n18342), .B(n18343), .X(n18341) );
  xor2_1 U17909 ( .A(n23995), .B(n12380), .X(n18343) );
  a21oi_1 U17910 ( .A1(n18182), .A2(n18344), .B1(n18183), .Y(n18342) );
  nand2_1 U17911 ( .A(n18345), .B(n12380), .Y(n18344) );
  xor2_1 U17912 ( .A(n18346), .B(n17915), .X(n18340) );
  inv_1 U17913 ( .A(n11523), .Y(n11715) );
  xor2_1 U17914 ( .A(n18347), .B(n18348), .X(n11523) );
  xor2_1 U17915 ( .A(n16832), .B(n18349), .X(n18348) );
  xor2_1 U17916 ( .A(n12968), .B(n12380), .X(n18349) );
  xor2_1 U17917 ( .A(n18350), .B(n18351), .X(n18347) );
  and2_0 U17918 ( .A(n18352), .B(n18353), .X(n18351) );
  xnor2_1 U17919 ( .A(n18163), .B(n18354), .Y(n11528) );
  xor2_1 U17920 ( .A(n12380), .B(n18355), .X(n18354) );
  a21oi_1 U17921 ( .A1(n18166), .A2(n18356), .B1(n18162), .Y(n18355) );
  o21ai_0 U17922 ( .A1(n12380), .A2(n18357), .B1(n18352), .Y(n18162) );
  xor2_1 U17923 ( .A(n18358), .B(n18359), .X(n18352) );
  nor2_1 U17924 ( .A(n18360), .B(n18183), .Y(n18359) );
  xor2_1 U17925 ( .A(n16914), .B(n18361), .X(n18183) );
  o21ai_0 U17926 ( .A1(n18192), .A2(n18193), .B1(n10826), .Y(n18361) );
  a21oi_1 U17927 ( .A1(n18346), .A2(n18362), .B1(n12380), .Y(n18360) );
  xor2_1 U17928 ( .A(n17644), .B(n18363), .X(n18357) );
  nor2_1 U17929 ( .A(n18356), .B(n18166), .Y(n18363) );
  inv_1 U17930 ( .A(n18353), .Y(n18356) );
  a21oi_1 U17931 ( .A1(n10826), .A2(n18182), .B1(n18165), .Y(n18353) );
  nor2_1 U17932 ( .A(n18179), .B(n18362), .Y(n18165) );
  inv_1 U17933 ( .A(n18178), .Y(n18362) );
  nand3_1 U17934 ( .A(n18192), .B(n18181), .C(n18182), .Y(n18179) );
  xor2_1 U17935 ( .A(n18364), .B(n17391), .X(n18182) );
  o21ai_0 U17936 ( .A1(n18193), .A2(n10826), .B1(n18339), .Y(n18364) );
  xor2_1 U17937 ( .A(n18365), .B(n12923), .X(n18339) );
  inv_1 U17938 ( .A(n16995), .Y(n12923) );
  o22ai_1 U17939 ( .A1(n18366), .A2(n18336), .B1(n12380), .B2(n18367), .Y(
        n18365) );
  nor2_1 U17940 ( .A(n18368), .B(n18335), .Y(n18367) );
  inv_1 U17941 ( .A(n18335), .Y(n18366) );
  nand2_1 U17942 ( .A(n18369), .B(n18331), .Y(n18335) );
  xnor2_1 U17943 ( .A(n18370), .B(n12806), .Y(n18331) );
  o211ai_1 U17944 ( .A1(n18328), .A2(n18371), .B1(n18372), .C1(n18373), .Y(
        n18370) );
  o21ai_0 U17945 ( .A1(n18329), .A2(n18374), .B1(n10607), .Y(n18372) );
  xor2_1 U17946 ( .A(n17031), .B(n18375), .X(n18369) );
  nand2_1 U17947 ( .A(n16015), .B(n18332), .Y(n18375) );
  o211ai_1 U17948 ( .A1(n18329), .A2(n18374), .B1(n18376), .C1(n18377), .Y(
        n18332) );
  o21ai_0 U17949 ( .A1(n18328), .A2(n18371), .B1(n23950), .Y(n18376) );
  inv_1 U17950 ( .A(n18328), .Y(n18374) );
  xor2_1 U17951 ( .A(n18378), .B(n18015), .X(n18328) );
  o21ai_0 U17952 ( .A1(n18379), .A2(n18324), .B1(n18322), .Y(n18378) );
  nand2_1 U17953 ( .A(n23938), .B(n18325), .Y(n18322) );
  xnor2_1 U17954 ( .A(n18380), .B(n10868), .Y(n18325) );
  inv_1 U17955 ( .A(n18379), .Y(n10868) );
  o211ai_1 U17956 ( .A1(n18319), .A2(n18320), .B1(n18381), .C1(n18382), .Y(
        n18380) );
  o21ai_0 U17957 ( .A1(n18383), .A2(n18384), .B1(n12320), .Y(n18381) );
  o211ai_1 U17958 ( .A1(n18383), .A2(n18384), .B1(n18385), .C1(n18386), .Y(
        n18324) );
  o21ai_0 U17959 ( .A1(n18319), .A2(n18320), .B1(n15953), .Y(n18385) );
  inv_1 U17960 ( .A(n18319), .Y(n18384) );
  xor2_1 U17961 ( .A(n18387), .B(n16850), .X(n18319) );
  o22ai_1 U17962 ( .A1(n18315), .A2(n18388), .B1(n23951), .B2(n18389), .Y(
        n18387) );
  nor2_1 U17963 ( .A(n18316), .B(n18390), .Y(n18389) );
  inv_1 U17964 ( .A(n18316), .Y(n18388) );
  xor2_1 U17965 ( .A(n18391), .B(n11048), .X(n18316) );
  o22ai_1 U17966 ( .A1(n18392), .A2(n18311), .B1(n18393), .B2(n15955), .Y(
        n18391) );
  nor2_1 U17967 ( .A(n18394), .B(n18312), .Y(n18393) );
  inv_1 U17968 ( .A(n18312), .Y(n18392) );
  o22ai_1 U17969 ( .A1(n18308), .A2(n18309), .B1(n23953), .B2(n18395), .Y(
        n18312) );
  and2_0 U17970 ( .A(n18309), .B(n18308), .X(n18395) );
  xor2_1 U17971 ( .A(n18396), .B(n18397), .X(n18308) );
  o22ai_1 U17972 ( .A1(n18398), .A2(n18303), .B1(n18399), .B2(n18305), .Y(
        n18396) );
  nor2_1 U17973 ( .A(n18400), .B(n18306), .Y(n18399) );
  inv_1 U17974 ( .A(n18306), .Y(n18398) );
  nand2_1 U17975 ( .A(n18401), .B(n18402), .Y(n18306) );
  xor2_1 U17976 ( .A(n18066), .B(n18403), .X(n18402) );
  nor2_1 U17977 ( .A(n18219), .B(n18221), .Y(n18403) );
  inv_1 U17978 ( .A(n18224), .Y(n18221) );
  o21ai_0 U17979 ( .A1(n12319), .A2(n18302), .B1(n18300), .Y(n18224) );
  xor2_1 U17980 ( .A(n18404), .B(n18405), .X(n18300) );
  nand2_1 U17981 ( .A(n18406), .B(n18407), .Y(n18404) );
  nor2_1 U17982 ( .A(n18407), .B(n18406), .Y(n18302) );
  nand2_1 U17983 ( .A(n18408), .B(n18231), .Y(n18407) );
  o211ai_1 U17984 ( .A1(n18298), .A2(n18409), .B1(n18410), .C1(n18411), .Y(
        n18231) );
  o21ai_0 U17985 ( .A1(n18296), .A2(n18412), .B1(n18413), .Y(n18410) );
  xor2_1 U17986 ( .A(n11413), .B(n18414), .X(n18408) );
  nand2_1 U17987 ( .A(n18230), .B(n16545), .Y(n18414) );
  xor2_1 U17988 ( .A(n18415), .B(n17774), .X(n18230) );
  o211ai_1 U17989 ( .A1(n18296), .A2(n18412), .B1(n18416), .C1(n18417), .Y(
        n18415) );
  o21ai_0 U17990 ( .A1(n18298), .A2(n18409), .B1(n23958), .Y(n18416) );
  inv_1 U17991 ( .A(n18412), .Y(n18298) );
  o22ai_1 U17992 ( .A1(n18293), .A2(n18295), .B1(n12393), .B2(n18418), .Y(
        n18412) );
  and2_0 U17993 ( .A(n18295), .B(n18293), .X(n18418) );
  o22ai_1 U17994 ( .A1(n18419), .A2(n18420), .B1(n1965), .B2(n18421), .Y(
        n18295) );
  nor2_1 U17995 ( .A(n18241), .B(n18240), .Y(n18421) );
  inv_1 U17996 ( .A(n18240), .Y(n18419) );
  o22ai_1 U17997 ( .A1(n18290), .A2(n18292), .B1(n12340), .B2(n18422), .Y(
        n18240) );
  and2_0 U17998 ( .A(n18292), .B(n18290), .X(n18422) );
  a21oi_1 U17999 ( .A1(n18287), .A2(n15990), .B1(n18423), .Y(n18290) );
  inv_1 U18000 ( .A(n18286), .Y(n18423) );
  xor2_1 U18001 ( .A(n12821), .B(n18424), .X(n18286) );
  nor2_1 U18002 ( .A(n18425), .B(n18426), .Y(n18424) );
  nand2_1 U18003 ( .A(n18425), .B(n18426), .Y(n18287) );
  a21oi_1 U18004 ( .A1(n18251), .A2(n23981), .B1(n18427), .Y(n18425) );
  inv_1 U18005 ( .A(n18250), .Y(n18427) );
  nand2_1 U18006 ( .A(n18428), .B(n18429), .Y(n18250) );
  xor2_1 U18007 ( .A(n16753), .B(n18430), .X(n18428) );
  nand2_1 U18008 ( .A(n18431), .B(n18432), .Y(n18251) );
  xor2_1 U18009 ( .A(n18430), .B(n17391), .X(n18431) );
  o22ai_1 U18010 ( .A1(n18283), .A2(n18433), .B1(n12394), .B2(n18434), .Y(
        n18430) );
  and2_0 U18011 ( .A(n18433), .B(n18283), .X(n18434) );
  inv_1 U18012 ( .A(n18284), .Y(n18433) );
  xor2_1 U18013 ( .A(n18435), .B(n11301), .X(n18283) );
  o22ai_1 U18014 ( .A1(n18257), .A2(n18256), .B1(n23987), .B2(n18436), .Y(
        n18435) );
  and2_0 U18015 ( .A(n18256), .B(n18257), .X(n18436) );
  a21oi_1 U18016 ( .A1(n18264), .A2(n23985), .B1(n18265), .Y(n18257) );
  xor2_1 U18017 ( .A(n17152), .B(n18437), .X(n18265) );
  nor2_1 U18018 ( .A(n18438), .B(n18439), .Y(n18437) );
  xnor2_1 U18019 ( .A(n18440), .B(n23995), .Y(n18264) );
  nand2_1 U18020 ( .A(n18438), .B(n18439), .Y(n18440) );
  a21oi_1 U18021 ( .A1(n15970), .A2(n18271), .B1(n18441), .Y(n18438) );
  inv_1 U18022 ( .A(n18270), .Y(n18441) );
  xor2_1 U18023 ( .A(n18442), .B(n18026), .X(n18270) );
  inv_1 U18024 ( .A(n16850), .Y(n18026) );
  nor3_1 U18025 ( .A(n13741), .B(n18443), .C(n18444), .Y(n16850) );
  nor2_1 U18026 ( .A(n18445), .B(n13956), .Y(n13741) );
  nand2_1 U18027 ( .A(n18446), .B(n18447), .Y(n18442) );
  xnor2_1 U18028 ( .A(n12956), .B(n18448), .Y(n18271) );
  nor2_1 U18029 ( .A(n18446), .B(n18447), .Y(n18448) );
  o22ai_1 U18030 ( .A1(n18449), .A2(n18450), .B1(n12305), .B2(n18281), .Y(
        n18447) );
  nor2_1 U18031 ( .A(n18279), .B(n16818), .Y(n18281) );
  inv_1 U18032 ( .A(n18449), .Y(n16818) );
  inv_1 U18033 ( .A(n18450), .Y(n18279) );
  xor2_1 U18034 ( .A(n18184), .B(n18451), .X(n18450) );
  a21oi_1 U18035 ( .A1(n18277), .A2(n18275), .B1(n18452), .Y(n18451) );
  inv_1 U18036 ( .A(n18276), .Y(n18452) );
  nand2_1 U18037 ( .A(n12401), .B(n16828), .Y(n18276) );
  inv_1 U18038 ( .A(n16824), .Y(n16828) );
  nand2_1 U18039 ( .A(n18453), .B(n18454), .Y(n18275) );
  nand3_1 U18040 ( .A(n18455), .B(n10608), .C(n17967), .Y(n18454) );
  xor2_1 U18041 ( .A(n17616), .B(n18456), .X(n18453) );
  nand2_1 U18042 ( .A(n18457), .B(n10775), .Y(n18456) );
  xor2_1 U18043 ( .A(n18458), .B(n18459), .X(n18457) );
  a21oi_1 U18044 ( .A1(n18460), .A2(n10608), .B1(n18461), .Y(n18459) );
  a21oi_1 U18045 ( .A1(n12331), .A2(n18462), .B1(n16842), .Y(n18461) );
  o21ai_0 U18046 ( .A1(n24022), .A2(n17966), .B1(n24019), .Y(n18460) );
  nand2_1 U18047 ( .A(n16824), .B(n18463), .Y(n18277) );
  xor2_1 U18048 ( .A(n18464), .B(n18465), .X(n16824) );
  xor2_1 U18049 ( .A(n11621), .B(n15895), .X(n18465) );
  nor2_1 U18050 ( .A(n18223), .B(n15931), .Y(n18219) );
  xor2_1 U18051 ( .A(n18466), .B(n18467), .X(n18401) );
  nand2_1 U18052 ( .A(n15931), .B(n18223), .Y(n18467) );
  o22ai_1 U18053 ( .A1(n13336), .A2(n13408), .B1(n18468), .B2(n13392), .Y(
        n17031) );
  nand2_1 U18054 ( .A(n11503), .B(n11703), .Y(n10819) );
  inv_1 U18055 ( .A(n10833), .Y(n11503) );
  nand2_1 U18056 ( .A(n18152), .B(n10832), .Y(n10833) );
  nand2_1 U18057 ( .A(n24052), .B(n12550), .Y(n10832) );
  nand2_1 U18058 ( .A(n24055), .B(n24052), .Y(n18152) );
  o21ai_0 U18059 ( .A1(n18469), .A2(n15459), .B1(inData[24]), .Y(n10821) );
  nor2_1 U18060 ( .A(n12550), .B(n11703), .Y(n15459) );
  nand2_1 U18061 ( .A(n12551), .B(n15863), .Y(n11703) );
  inv_1 U18062 ( .A(n24052), .Y(n12551) );
  inv_1 U18063 ( .A(n11177), .Y(n18469) );
  nand2_1 U18064 ( .A(n11618), .B(n24052), .Y(n11177) );
  inv_1 U18065 ( .A(n11226), .Y(n11618) );
  nand2_1 U18066 ( .A(n15863), .B(n12550), .Y(n11226) );
  inv_1 U18067 ( .A(n24062), .Y(n12550) );
  inv_1 U18068 ( .A(n24055), .Y(n15863) );
  nor2_1 U18069 ( .A(n10774), .B(n18470), .Y(n10145) );
  xor2_1 U18070 ( .A(n12951), .B(n18471), .X(n18470) );
  nand2_1 U18071 ( .A(n12950), .B(n12948), .Y(n18471) );
  nand2_1 U18072 ( .A(n18472), .B(n18473), .Y(n12948) );
  xor2_1 U18073 ( .A(n18474), .B(n16742), .X(n12950) );
  nand2_1 U18074 ( .A(n18475), .B(n18476), .Y(n18474) );
  xor2_1 U18075 ( .A(n18472), .B(n18477), .X(n18475) );
  xnor2_1 U18076 ( .A(n18478), .B(n12961), .Y(n18472) );
  mux2i_1 U18077 ( .A0(n18479), .A1(n18480), .S(n18077), .Y(n12961) );
  o22ai_1 U18078 ( .A1(n23949), .A2(n18481), .B1(n811), .B2(n18482), .Y(n18480) );
  nor2_1 U18079 ( .A(n16015), .B(n18483), .Y(n18482) );
  nand2_1 U18080 ( .A(n18484), .B(n18483), .Y(n18479) );
  xor2_1 U18081 ( .A(n12429), .B(n10826), .X(n18478) );
  o22ai_1 U18082 ( .A1(n11410), .A2(n11409), .B1(n18485), .B2(n11411), .Y(
        n12951) );
  and2_0 U18083 ( .A(n11409), .B(n11410), .X(n18485) );
  o22ai_1 U18084 ( .A1(n18486), .A2(n18487), .B1(n18488), .B2(n12940), .Y(
        n11409) );
  nand2_1 U18085 ( .A(n18489), .B(n12971), .Y(n12940) );
  nand2_1 U18086 ( .A(n18490), .B(n18491), .Y(n12971) );
  xor2_1 U18087 ( .A(n16666), .B(n18492), .X(n18489) );
  nand2_1 U18088 ( .A(n12966), .B(n18493), .Y(n18492) );
  inv_1 U18089 ( .A(n12973), .Y(n18493) );
  nor2_1 U18090 ( .A(n18490), .B(n18491), .Y(n12973) );
  xnor2_1 U18091 ( .A(n18494), .B(n18495), .Y(n18490) );
  xor2_1 U18092 ( .A(n18496), .B(n16493), .X(n12966) );
  o22ai_1 U18093 ( .A1(n11467), .A2(n11465), .B1(n11464), .B2(n18497), .Y(
        n18496) );
  and2_0 U18094 ( .A(n18498), .B(n11467), .X(n18497) );
  a21oi_1 U18095 ( .A1(n18499), .A2(n17233), .B1(n17234), .Y(n11464) );
  and2_0 U18096 ( .A(n18500), .B(n18501), .X(n17234) );
  inv_1 U18097 ( .A(n18502), .Y(n17233) );
  o22ai_1 U18098 ( .A1(n17044), .A2(n17046), .B1(n18503), .B2(n17047), .Y(
        n18502) );
  and2_0 U18099 ( .A(n17046), .B(n17044), .X(n18503) );
  o22ai_1 U18100 ( .A1(n17040), .A2(n17042), .B1(n18504), .B2(n17041), .Y(
        n17046) );
  inv_1 U18101 ( .A(n18505), .Y(n17041) );
  and2_0 U18102 ( .A(n17042), .B(n17040), .X(n18504) );
  o22ai_1 U18103 ( .A1(n11220), .A2(n11222), .B1(n18506), .B2(n11223), .Y(
        n17042) );
  and2_0 U18104 ( .A(n11222), .B(n11220), .X(n18506) );
  o22ai_1 U18105 ( .A1(n12538), .A2(n12539), .B1(n18507), .B2(n18508), .Y(
        n11222) );
  and2_0 U18106 ( .A(n12539), .B(n12538), .X(n18507) );
  o22ai_1 U18107 ( .A1(n18509), .A2(n18510), .B1(n18511), .B2(n18512), .Y(
        n12539) );
  and2_0 U18108 ( .A(n18513), .B(n18514), .X(n18511) );
  a21oi_1 U18109 ( .A1(n11275), .A2(n11274), .B1(n18515), .Y(n12538) );
  inv_1 U18110 ( .A(n11276), .Y(n18515) );
  nand2_1 U18111 ( .A(n18516), .B(n18517), .Y(n11276) );
  xnor2_1 U18112 ( .A(n16275), .B(n18518), .Y(n18516) );
  mux2_1 U18113 ( .A0(n18519), .A1(n18520), .S(n18521), .X(n11274) );
  nand2_1 U18114 ( .A(n17034), .B(n18522), .Y(n18520) );
  and2_0 U18115 ( .A(n18523), .B(n18524), .X(n17034) );
  o21ai_0 U18116 ( .A1(n17458), .A2(n18525), .B1(n18526), .Y(n18524) );
  o221ai_1 U18117 ( .A1(n18527), .A2(n18525), .B1(n17037), .B2(n18526), .C1(
        n18523), .Y(n18519) );
  or3_1 U18118 ( .A(n18526), .B(n17458), .C(n18525), .X(n18523) );
  inv_1 U18119 ( .A(n18522), .Y(n17037) );
  a21oi_1 U18120 ( .A1(n18526), .A2(n17458), .B1(n18522), .Y(n18527) );
  o21ai_0 U18121 ( .A1(n11163), .A2(n18528), .B1(n18529), .Y(n18522) );
  xor2_1 U18122 ( .A(n14685), .B(n18530), .X(n18529) );
  nand2_1 U18123 ( .A(n11165), .B(n11167), .Y(n18530) );
  nand2_1 U18124 ( .A(n18531), .B(n18528), .Y(n11167) );
  xor2_1 U18125 ( .A(n18532), .B(n11166), .X(n18531) );
  o21ai_0 U18126 ( .A1(n18533), .A2(n11300), .B1(n11302), .Y(n11165) );
  xor2_1 U18127 ( .A(n18534), .B(n18535), .X(n11302) );
  or2_0 U18128 ( .A(n18536), .B(n18537), .X(n18534) );
  o22ai_1 U18129 ( .A1(n12495), .A2(n18538), .B1(n18539), .B2(n12497), .Y(
        n11300) );
  o22ai_1 U18130 ( .A1(n12527), .A2(n12528), .B1(n18540), .B2(n18541), .Y(
        n12497) );
  and2_0 U18131 ( .A(n12528), .B(n12527), .X(n18540) );
  xnor2_1 U18132 ( .A(n18542), .B(n18543), .Y(n12528) );
  xor2_1 U18133 ( .A(n17133), .B(n18544), .X(n18542) );
  a21oi_1 U18134 ( .A1(n12340), .A2(n11149), .B1(n18545), .Y(n18544) );
  xor2_1 U18135 ( .A(n18546), .B(n18052), .X(n12527) );
  o22ai_1 U18136 ( .A1(n18547), .A2(n12483), .B1(n12489), .B2(n18548), .Y(
        n18546) );
  nor2_1 U18137 ( .A(n18549), .B(n12488), .Y(n18548) );
  inv_1 U18138 ( .A(n12483), .Y(n18549) );
  xor2_1 U18139 ( .A(n18550), .B(n18551), .X(n12483) );
  xor2_1 U18140 ( .A(n12392), .B(n12376), .X(n18551) );
  xor2_1 U18141 ( .A(n11428), .B(n18552), .X(n18550) );
  inv_1 U18142 ( .A(n12488), .Y(n18547) );
  o21ai_0 U18143 ( .A1(n12824), .A2(n18553), .B1(n12820), .Y(n12488) );
  nand2_1 U18144 ( .A(n18554), .B(n18555), .Y(n12820) );
  xor2_1 U18145 ( .A(n23979), .B(n12822), .X(n18553) );
  nor2_1 U18146 ( .A(n18554), .B(n18555), .Y(n12822) );
  xnor2_1 U18147 ( .A(n18556), .B(n18557), .Y(n18554) );
  a21oi_1 U18148 ( .A1(n11354), .A2(n11350), .B1(n11353), .Y(n12824) );
  xor2_1 U18149 ( .A(n18521), .B(n18558), .X(n11353) );
  nor2_1 U18150 ( .A(n18559), .B(n18560), .Y(n18558) );
  inv_1 U18151 ( .A(n18561), .Y(n11350) );
  a21oi_1 U18152 ( .A1(n11555), .A2(n11557), .B1(n18562), .Y(n18561) );
  inv_1 U18153 ( .A(n11556), .Y(n18562) );
  xor2_1 U18154 ( .A(n18563), .B(n18564), .X(n11556) );
  nor2_1 U18155 ( .A(n18565), .B(n18566), .Y(n18564) );
  nand2_1 U18156 ( .A(n18567), .B(n18566), .Y(n11557) );
  xnor2_1 U18157 ( .A(n18568), .B(n18569), .Y(n18566) );
  nor2_1 U18158 ( .A(n18570), .B(n18571), .Y(n18569) );
  xor2_1 U18159 ( .A(n11159), .B(n18565), .X(n18567) );
  o21ai_0 U18160 ( .A1(n18572), .A2(n11575), .B1(n11577), .Y(n11555) );
  xnor2_1 U18161 ( .A(n16801), .B(n18573), .Y(n11577) );
  nor2_1 U18162 ( .A(n18574), .B(n18575), .Y(n18573) );
  inv_1 U18163 ( .A(n18576), .Y(n18574) );
  o22ai_1 U18164 ( .A1(n12790), .A2(n12787), .B1(n18577), .B2(n12789), .Y(
        n11575) );
  and2_0 U18165 ( .A(n12787), .B(n12790), .X(n18577) );
  mux2_1 U18166 ( .A0(n18578), .A1(n18579), .S(n11428), .X(n12787) );
  nand2_1 U18167 ( .A(n18580), .B(n17029), .Y(n18579) );
  xnor2_1 U18168 ( .A(n18581), .B(n18582), .Y(n17029) );
  o22ai_1 U18169 ( .A1(n18583), .A2(n17032), .B1(n18584), .B2(n18581), .Y(
        n18578) );
  xor2_1 U18170 ( .A(n18585), .B(n18586), .X(n18581) );
  xor2_1 U18171 ( .A(n18587), .B(n18588), .X(n18586) );
  xor2_1 U18172 ( .A(n18589), .B(n11710), .X(n18585) );
  nor2_1 U18173 ( .A(n18580), .B(n18582), .Y(n18584) );
  inv_1 U18174 ( .A(n17032), .Y(n18580) );
  o22ai_1 U18175 ( .A1(n17239), .A2(n17241), .B1(n18590), .B2(n17237), .Y(
        n17032) );
  o21ai_0 U18176 ( .A1(n12810), .A2(n12813), .B1(n12811), .Y(n17237) );
  xnor2_1 U18177 ( .A(n18591), .B(n16931), .Y(n12811) );
  nand2_1 U18178 ( .A(n18592), .B(n18593), .Y(n18591) );
  xor2_1 U18179 ( .A(n10919), .B(n18594), .X(n12813) );
  nor2_1 U18180 ( .A(n18592), .B(n18593), .Y(n18594) );
  xor2_1 U18181 ( .A(n18595), .B(n23993), .X(n18592) );
  nand2_1 U18182 ( .A(n18596), .B(n18597), .Y(n18595) );
  a21oi_1 U18183 ( .A1(n11784), .A2(n11782), .B1(n18598), .Y(n12810) );
  inv_1 U18184 ( .A(n11783), .Y(n18598) );
  xor2_1 U18185 ( .A(n18021), .B(n18599), .X(n11783) );
  nor2_1 U18186 ( .A(n18600), .B(n18601), .Y(n18599) );
  and3_1 U18187 ( .A(n18602), .B(n18603), .C(n18604), .X(n11782) );
  nor3_1 U18188 ( .A(n18605), .B(n18606), .C(n18607), .Y(n18604) );
  xor2_1 U18189 ( .A(n13401), .B(n18608), .X(n18603) );
  nand2_1 U18190 ( .A(n18609), .B(n12464), .Y(n18608) );
  xor2_1 U18191 ( .A(n17458), .B(n18610), .X(n18602) );
  and2_0 U18192 ( .A(n12506), .B(n18611), .X(n18610) );
  nand2_1 U18193 ( .A(n18600), .B(n18601), .Y(n11784) );
  xor2_1 U18194 ( .A(n18612), .B(n10608), .X(n18601) );
  o21ai_0 U18195 ( .A1(n10639), .A2(n18613), .B1(n18614), .Y(n18612) );
  and2_0 U18196 ( .A(n17241), .B(n18615), .X(n18590) );
  xnor2_1 U18197 ( .A(n18616), .B(n18617), .Y(n17241) );
  nand2_1 U18198 ( .A(n18618), .B(n18619), .Y(n18616) );
  inv_1 U18199 ( .A(n18620), .Y(n18618) );
  xor2_1 U18200 ( .A(n18615), .B(n12881), .X(n17239) );
  xor2_1 U18201 ( .A(n18621), .B(n18622), .X(n12790) );
  xor2_1 U18202 ( .A(n12549), .B(n12388), .X(n18622) );
  xor2_1 U18203 ( .A(n18623), .B(n18624), .X(n18621) );
  xor2_1 U18204 ( .A(n12297), .B(n11578), .X(n18572) );
  nand2_1 U18205 ( .A(n18625), .B(n18575), .Y(n11578) );
  xnor2_1 U18206 ( .A(n18626), .B(n18627), .Y(n18575) );
  xor2_1 U18207 ( .A(n23985), .B(n12547), .X(n18627) );
  xnor2_1 U18208 ( .A(n18628), .B(n12686), .Y(n18626) );
  xor2_1 U18209 ( .A(n18576), .B(n17715), .X(n18625) );
  nand2_1 U18210 ( .A(n18560), .B(n18559), .Y(n11354) );
  xor2_1 U18211 ( .A(n18629), .B(n18630), .X(n18560) );
  xor2_1 U18212 ( .A(n10631), .B(n12394), .X(n18629) );
  nor2_1 U18213 ( .A(n12496), .B(n18631), .Y(n18539) );
  inv_1 U18214 ( .A(n12495), .Y(n18631) );
  inv_1 U18215 ( .A(n18538), .Y(n12496) );
  xor2_1 U18216 ( .A(n18632), .B(n18633), .X(n18538) );
  xor2_1 U18217 ( .A(n16845), .B(n18634), .X(n18633) );
  xor2_1 U18218 ( .A(n23932), .B(n10606), .X(n18632) );
  xor2_1 U18219 ( .A(n18635), .B(n11048), .X(n12495) );
  inv_1 U18220 ( .A(n11303), .Y(n18533) );
  nand2_1 U18221 ( .A(n18636), .B(n18536), .Y(n11303) );
  xnor2_1 U18222 ( .A(n18637), .B(n18638), .Y(n18536) );
  nor2_1 U18223 ( .A(n18639), .B(n18640), .Y(n18638) );
  inv_1 U18224 ( .A(n18641), .Y(n18639) );
  xor2_1 U18225 ( .A(n18642), .B(n17915), .X(n18636) );
  inv_1 U18226 ( .A(n11164), .Y(n18528) );
  xor2_1 U18227 ( .A(n18643), .B(n18644), .X(n11164) );
  xor2_1 U18228 ( .A(n18645), .B(n24045), .X(n18643) );
  xor2_1 U18229 ( .A(n18646), .B(n18647), .X(n18526) );
  xor2_1 U18230 ( .A(n23959), .B(n12373), .X(n18647) );
  nand2_1 U18231 ( .A(n18648), .B(n18518), .Y(n11275) );
  xnor2_1 U18232 ( .A(n18649), .B(n18650), .Y(n18518) );
  xor2_1 U18233 ( .A(n63), .B(n12319), .X(n18650) );
  xor2_1 U18234 ( .A(n18651), .B(n18517), .X(n18648) );
  inv_1 U18235 ( .A(n18652), .Y(n18517) );
  xnor2_1 U18236 ( .A(n18653), .B(n18654), .Y(n11220) );
  xor2_1 U18237 ( .A(n67), .B(n23948), .X(n18654) );
  xor2_1 U18238 ( .A(n18655), .B(n18656), .X(n17040) );
  xnor2_1 U18239 ( .A(n18657), .B(n18658), .Y(n17044) );
  nand2_1 U18240 ( .A(n18659), .B(n18660), .Y(n18657) );
  inv_1 U18241 ( .A(n18661), .Y(n18660) );
  inv_1 U18242 ( .A(n17235), .Y(n18499) );
  xor2_1 U18243 ( .A(n17644), .B(n18662), .X(n17235) );
  nor2_1 U18244 ( .A(n18501), .B(n18500), .Y(n18662) );
  xor2_1 U18245 ( .A(n18663), .B(n18664), .X(n18500) );
  nand2_1 U18246 ( .A(n18665), .B(n18666), .Y(n18663) );
  inv_1 U18247 ( .A(n18667), .Y(n18665) );
  o211ai_1 U18248 ( .A1(n18668), .A2(n18445), .B1(n13764), .C1(n16146), .Y(
        n17644) );
  xor2_1 U18249 ( .A(n11466), .B(n12297), .X(n11465) );
  xor2_1 U18250 ( .A(n18669), .B(n18670), .X(n11467) );
  nor2_1 U18251 ( .A(n12938), .B(n18671), .Y(n18488) );
  xor2_1 U18252 ( .A(n12939), .B(n12936), .X(n18671) );
  inv_1 U18253 ( .A(n18015), .Y(n12939) );
  a211oi_1 U18254 ( .A1(n24013), .A2(n18672), .B1(n13275), .C1(n18673), .Y(
        n18015) );
  nor2_1 U18255 ( .A(n13408), .B(n13403), .Y(n13275) );
  inv_1 U18256 ( .A(n12936), .Y(n18487) );
  xor2_1 U18257 ( .A(n18674), .B(n18675), .X(n12936) );
  xor2_1 U18258 ( .A(n18676), .B(n18677), .X(n18675) );
  nand2_1 U18259 ( .A(n18678), .B(n18679), .Y(n18676) );
  xor2_1 U18260 ( .A(n18680), .B(n12297), .X(n18674) );
  xor2_1 U18261 ( .A(n18484), .B(n18481), .X(n11410) );
  inv_1 U18262 ( .A(n18483), .Y(n18481) );
  o21ai_0 U18263 ( .A1(n18681), .A2(n18677), .B1(n18678), .Y(n18483) );
  xor2_1 U18264 ( .A(n18682), .B(n18683), .X(n18678) );
  nor2_1 U18265 ( .A(n10607), .B(n16959), .Y(n18683) );
  mux2i_1 U18266 ( .A0(n18684), .A1(n18685), .S(n17475), .Y(n18677) );
  o22ai_1 U18267 ( .A1(n23938), .A2(n18494), .B1(n68), .B2(n18686), .Y(n18685)
         );
  nor2_1 U18268 ( .A(n16013), .B(n18687), .Y(n18686) );
  nand2_1 U18269 ( .A(n18687), .B(n18495), .Y(n18684) );
  xnor2_1 U18270 ( .A(n68), .B(n16013), .Y(n18495) );
  inv_1 U18271 ( .A(n18494), .Y(n18687) );
  mux2i_1 U18272 ( .A0(n18688), .A1(n18689), .S(n17830), .Y(n18494) );
  nand2_1 U18273 ( .A(n18669), .B(n18690), .Y(n18689) );
  xor2_1 U18274 ( .A(n16966), .B(n12320), .X(n18669) );
  o22ai_1 U18275 ( .A1(n12320), .A2(n18670), .B1(n18691), .B2(n16966), .Y(
        n18688) );
  inv_1 U18276 ( .A(n23920), .Y(n16966) );
  nor2_1 U18277 ( .A(n15953), .B(n18690), .Y(n18691) );
  inv_1 U18278 ( .A(n18690), .Y(n18670) );
  o21ai_0 U18279 ( .A1(n18664), .A2(n18667), .B1(n18666), .Y(n18690) );
  nand2_1 U18280 ( .A(n23951), .B(n18692), .Y(n18666) );
  xor2_1 U18281 ( .A(n11574), .B(n18693), .X(n18667) );
  nor2_1 U18282 ( .A(n23951), .B(n18692), .Y(n18693) );
  inv_1 U18283 ( .A(n64), .Y(n18692) );
  a21oi_1 U18284 ( .A1(n18659), .A2(n18658), .B1(n18661), .Y(n18664) );
  nor2_1 U18285 ( .A(n15955), .B(n4), .Y(n18661) );
  mux2_1 U18286 ( .A0(n18694), .A1(n18695), .S(n17620), .X(n18658) );
  nand2_1 U18287 ( .A(n18696), .B(n18656), .Y(n18695) );
  xor2_1 U18288 ( .A(n771), .B(n23953), .X(n18656) );
  o22ai_1 U18289 ( .A1(n23953), .A2(n18655), .B1(n771), .B2(n18697), .Y(n18694) );
  nor2_1 U18290 ( .A(n18696), .B(n16611), .Y(n18697) );
  inv_1 U18291 ( .A(n18655), .Y(n18696) );
  o22ai_1 U18292 ( .A1(n23948), .A2(n18698), .B1(n67), .B2(n18699), .Y(n18655)
         );
  nor2_1 U18293 ( .A(n18653), .B(n18305), .Y(n18699) );
  inv_1 U18294 ( .A(n18653), .Y(n18698) );
  xor2_1 U18295 ( .A(n18700), .B(n11103), .X(n18653) );
  nand2_1 U18296 ( .A(n18513), .B(n18510), .Y(n18700) );
  nand2_1 U18297 ( .A(n18514), .B(n18512), .Y(n18510) );
  o22ai_1 U18298 ( .A1(n12319), .A2(n18649), .B1(n18701), .B2(n18702), .Y(
        n18512) );
  inv_1 U18299 ( .A(n63), .Y(n18702) );
  and2_0 U18300 ( .A(n12319), .B(n18649), .X(n18701) );
  xor2_1 U18301 ( .A(n18703), .B(n23903), .X(n18649) );
  o22ai_1 U18302 ( .A1(n18704), .A2(n11212), .B1(n23959), .B2(n18705), .Y(
        n18703) );
  nor2_1 U18303 ( .A(n12373), .B(n18646), .Y(n18705) );
  inv_1 U18304 ( .A(n12373), .Y(n11212) );
  inv_1 U18305 ( .A(n18646), .Y(n18704) );
  xor2_1 U18306 ( .A(n12968), .B(n18706), .X(n18646) );
  mux2i_1 U18307 ( .A0(n18707), .A1(n18708), .S(n10928), .Y(n18706) );
  and2_0 U18308 ( .A(n18709), .B(n18644), .X(n18708) );
  xor2_1 U18309 ( .A(n11288), .B(n18413), .X(n18644) );
  o22ai_1 U18310 ( .A1(n12511), .A2(n18709), .B1(n23958), .B2(n18710), .Y(
        n18707) );
  nor2_1 U18311 ( .A(n18645), .B(n11288), .Y(n18710) );
  inv_1 U18312 ( .A(n12511), .Y(n11288) );
  inv_1 U18313 ( .A(n18645), .Y(n18709) );
  xor2_1 U18314 ( .A(n11601), .B(n18711), .X(n18645) );
  a21oi_1 U18315 ( .A1(n18637), .A2(n18641), .B1(n18640), .Y(n18711) );
  xor2_1 U18316 ( .A(n16464), .B(n18712), .X(n18640) );
  nor2_1 U18317 ( .A(n62), .B(n15902), .Y(n18712) );
  nand2_1 U18318 ( .A(n62), .B(n15902), .Y(n18641) );
  o22ai_1 U18319 ( .A1(n1965), .A2(n18634), .B1(n23932), .B2(n18713), .Y(
        n18637) );
  and2_0 U18320 ( .A(n18634), .B(n1965), .X(n18713) );
  o32ai_1 U18321 ( .A1(n18034), .A2(n23928), .A3(n16510), .B1(n18543), .B2(
        n18545), .Y(n18634) );
  xor2_1 U18322 ( .A(n18034), .B(n18714), .X(n18545) );
  nor2_1 U18323 ( .A(n12340), .B(n11149), .Y(n18714) );
  inv_1 U18324 ( .A(n23928), .Y(n11149) );
  inv_1 U18325 ( .A(n18715), .Y(n18543) );
  o22ai_1 U18326 ( .A1(n12376), .A2(n18552), .B1(n18716), .B2(n15990), .Y(
        n18715) );
  nor2_1 U18327 ( .A(n18717), .B(n12746), .Y(n18716) );
  inv_1 U18328 ( .A(n12376), .Y(n12746) );
  inv_1 U18329 ( .A(n18717), .Y(n18552) );
  mux2i_1 U18330 ( .A0(n18718), .A1(n18719), .S(n17952), .Y(n18717) );
  inv_1 U18331 ( .A(n11668), .Y(n17952) );
  o22ai_1 U18332 ( .A1(n18557), .A2(n15999), .B1(n53), .B2(n18720), .Y(n18719)
         );
  nor2_1 U18333 ( .A(n23981), .B(n18721), .Y(n18720) );
  inv_1 U18334 ( .A(n18721), .Y(n18557) );
  nand2_1 U18335 ( .A(n18556), .B(n18721), .Y(n18718) );
  o22ai_1 U18336 ( .A1(n12394), .A2(n18630), .B1(n18722), .B2(n10631), .Y(
        n18721) );
  and2_0 U18337 ( .A(n12394), .B(n18630), .X(n18722) );
  a21oi_1 U18338 ( .A1(n18723), .A2(n18568), .B1(n18571), .Y(n18630) );
  xnor2_1 U18339 ( .A(n18724), .B(n18725), .Y(n18571) );
  and2_0 U18340 ( .A(n16453), .B(n12520), .X(n18725) );
  o22ai_1 U18341 ( .A1(n18628), .A2(n17017), .B1(n18726), .B2(n18262), .Y(
        n18568) );
  and2_0 U18342 ( .A(n18628), .B(n17017), .X(n18726) );
  inv_1 U18343 ( .A(n12547), .Y(n17017) );
  o22ai_1 U18344 ( .A1(n18623), .A2(n15970), .B1(n12549), .B2(n18727), .Y(
        n18628) );
  and2_0 U18345 ( .A(n15970), .B(n18623), .X(n18727) );
  mux2i_1 U18346 ( .A0(n18728), .A1(n18729), .S(n16902), .Y(n18623) );
  o22ai_1 U18347 ( .A1(n15972), .A2(n18730), .B1(n49), .B2(n18731), .Y(n18729)
         );
  nor2_1 U18348 ( .A(n12305), .B(n18589), .Y(n18731) );
  inv_1 U18349 ( .A(n18589), .Y(n18730) );
  nor2_1 U18350 ( .A(n18587), .B(n18589), .Y(n18728) );
  xor2_1 U18351 ( .A(n18732), .B(n18733), .X(n18589) );
  a21oi_1 U18352 ( .A1(n18617), .A2(n18619), .B1(n18620), .Y(n18733) );
  xor2_1 U18353 ( .A(n18734), .B(n18052), .X(n18620) );
  nand2_1 U18354 ( .A(n46), .B(n12401), .Y(n18734) );
  or2_0 U18355 ( .A(n46), .B(n12401), .X(n18619) );
  a21oi_1 U18356 ( .A1(n18596), .A2(n23993), .B1(n18735), .Y(n18617) );
  inv_1 U18357 ( .A(n18597), .Y(n18735) );
  nand2_1 U18358 ( .A(n58), .B(n18736), .Y(n18597) );
  nand3_1 U18359 ( .A(n15916), .B(n18614), .C(n18737), .Y(n18736) );
  nand4_1 U18360 ( .A(n18737), .B(n15916), .C(n18614), .D(n11776), .Y(n18596)
         );
  inv_1 U18361 ( .A(n58), .Y(n11776) );
  nand2_1 U18362 ( .A(n18613), .B(n10639), .Y(n18614) );
  nand2_1 U18363 ( .A(n18738), .B(n15913), .Y(n18613) );
  nand2_1 U18364 ( .A(n24011), .B(n24022), .Y(n15916) );
  inv_1 U18365 ( .A(n18739), .Y(n18737) );
  a21oi_1 U18366 ( .A1(n18738), .A2(n821), .B1(n10608), .Y(n18739) );
  xor2_1 U18367 ( .A(n49), .B(n12305), .X(n18587) );
  inv_1 U18368 ( .A(n18570), .Y(n18723) );
  nor2_1 U18369 ( .A(n16453), .B(n12520), .Y(n18570) );
  xor2_1 U18370 ( .A(n53), .B(n15999), .X(n18556) );
  xnor2_1 U18371 ( .A(n11574), .B(n18740), .Y(n18514) );
  and2_0 U18372 ( .A(n12302), .B(n12484), .X(n18740) );
  inv_1 U18373 ( .A(n18509), .Y(n18513) );
  nor2_1 U18374 ( .A(n12302), .B(n12484), .Y(n18509) );
  xnor2_1 U18375 ( .A(n18680), .B(n18741), .Y(n18659) );
  and2_0 U18376 ( .A(n15955), .B(n4), .X(n18741) );
  inv_1 U18377 ( .A(n18679), .Y(n18681) );
  nand2_1 U18378 ( .A(n10607), .B(n16959), .Y(n18679) );
  inv_1 U18379 ( .A(n12580), .Y(n16959) );
  xor2_1 U18380 ( .A(n811), .B(n23949), .X(n18484) );
  inv_1 U18381 ( .A(n23922), .Y(n10774) );
  nand2_1 U18382 ( .A(n18742), .B(n15877), .Y(n10144) );
  nand3_1 U18383 ( .A(n11482), .B(n11150), .C(n24054), .Y(n15877) );
  mux2i_1 U18384 ( .A0(n18743), .A1(n18744), .S(n11482), .Y(n18742) );
  xor2_1 U18385 ( .A(n18745), .B(n18746), .X(n18744) );
  xor2_1 U18386 ( .A(n811), .B(n779), .X(n18746) );
  nand2_1 U18387 ( .A(n12429), .B(n11679), .Y(n18745) );
  inv_1 U18388 ( .A(n12467), .Y(n11679) );
  xor2_1 U18389 ( .A(n18747), .B(n18748), .X(n18743) );
  xnor2_1 U18390 ( .A(n23997), .B(n16739), .Y(n18748) );
  nand3_1 U18391 ( .A(n18749), .B(n18750), .C(n23922), .Y(n10143) );
  o21ai_0 U18392 ( .A1(n10953), .A2(n10954), .B1(n18751), .Y(n18750) );
  inv_1 U18393 ( .A(n10956), .Y(n18751) );
  o211ai_1 U18394 ( .A1(n18458), .A2(n10953), .B1(n18752), .C1(n18753), .Y(
        n10956) );
  o21ai_0 U18395 ( .A1(n18754), .A2(n18755), .B1(n18756), .Y(n18749) );
  inv_1 U18396 ( .A(n18752), .Y(n18756) );
  o22ai_1 U18397 ( .A1(n18757), .A2(n18758), .B1(n18759), .B2(n18760), .Y(
        n18752) );
  and2_0 U18398 ( .A(n18758), .B(n18757), .X(n18759) );
  inv_1 U18399 ( .A(n18753), .Y(n18755) );
  nand3_1 U18400 ( .A(n18458), .B(n10954), .C(n10953), .Y(n18753) );
  a21oi_1 U18401 ( .A1(n18458), .A2(n10954), .B1(n10953), .Y(n18754) );
  xor2_1 U18402 ( .A(n18761), .B(n10813), .X(n10953) );
  inv_1 U18403 ( .A(n10810), .Y(n10813) );
  xor2_1 U18404 ( .A(n17573), .B(n18762), .X(n10810) );
  a21oi_1 U18405 ( .A1(n18763), .A2(n18764), .B1(n18765), .Y(n18762) );
  xnor2_1 U18406 ( .A(n10951), .B(n3), .Y(n18761) );
  a21oi_1 U18407 ( .A1(n18766), .A2(n18767), .B1(n18768), .Y(n10951) );
  o21ai_0 U18408 ( .A1(n18769), .A2(n10948), .B1(n18770), .Y(n10954) );
  mux2i_1 U18409 ( .A0(n10944), .A1(n18771), .S(n10945), .Y(n18770) );
  nor2_1 U18410 ( .A(n10970), .B(n10949), .Y(n18771) );
  nor2_1 U18411 ( .A(n10884), .B(n10970), .Y(n10944) );
  xor2_1 U18412 ( .A(n10945), .B(n10949), .X(n18769) );
  inv_1 U18413 ( .A(n10884), .Y(n10949) );
  xor2_1 U18414 ( .A(n18772), .B(n18773), .X(n10884) );
  xor2_1 U18415 ( .A(n11520), .B(n10938), .X(n18773) );
  o21ai_0 U18416 ( .A1(outData[31]), .A2(n18774), .B1(n18775), .Y(n10938) );
  xor2_1 U18417 ( .A(n11428), .B(n18776), .X(n18775) );
  nand2_1 U18418 ( .A(n18777), .B(n18778), .Y(n18776) );
  inv_1 U18419 ( .A(n10840), .Y(n11428) );
  nand2_1 U18420 ( .A(n10937), .B(n10939), .Y(n18772) );
  nand2_1 U18421 ( .A(n18779), .B(n18124), .Y(n10939) );
  xor2_1 U18422 ( .A(n17475), .B(n18780), .X(n10937) );
  nor2_1 U18423 ( .A(n18124), .B(n18779), .Y(n18780) );
  o22ai_1 U18424 ( .A1(n18781), .A2(n10948), .B1(n18782), .B2(n18783), .Y(
        n10945) );
  nor2_1 U18425 ( .A(n18784), .B(n10970), .Y(n18782) );
  inv_1 U18426 ( .A(n10948), .Y(n10970) );
  nand2_1 U18427 ( .A(n23922), .B(n18785), .Y(n10142) );
  xnor2_1 U18428 ( .A(n18760), .B(n18786), .Y(n18785) );
  xor2_1 U18429 ( .A(n18757), .B(n18758), .X(n18786) );
  xnor2_1 U18430 ( .A(n18787), .B(n18783), .Y(n18758) );
  xor2_1 U18431 ( .A(n10948), .B(n18784), .X(n18787) );
  inv_1 U18432 ( .A(n18781), .Y(n18784) );
  o21ai_0 U18433 ( .A1(n18788), .A2(n18789), .B1(n18790), .Y(n18781) );
  xor2_1 U18434 ( .A(n17573), .B(n18791), .X(n18790) );
  nand2_1 U18435 ( .A(n11697), .B(n18792), .Y(n18791) );
  nor2_1 U18436 ( .A(n11697), .B(n18792), .Y(n18789) );
  o21ai_0 U18437 ( .A1(outData[31]), .A2(n18793), .B1(n18794), .Y(n10948) );
  mux2i_1 U18438 ( .A0(n18795), .A1(n18796), .S(n18777), .Y(n18794) );
  nor2_1 U18439 ( .A(n18774), .B(n18124), .Y(n18796) );
  inv_1 U18440 ( .A(n18778), .Y(n18795) );
  nand2_1 U18441 ( .A(outData[31]), .B(n18774), .Y(n18778) );
  xor2_1 U18442 ( .A(n18777), .B(n18774), .X(n18793) );
  o22ai_1 U18443 ( .A1(n18797), .A2(n18798), .B1(outData[31]), .B2(n18799), 
        .Y(n18777) );
  nor2_1 U18444 ( .A(n18800), .B(n18801), .Y(n18799) );
  xor2_1 U18445 ( .A(n14685), .B(n18802), .X(n18757) );
  a21oi_1 U18446 ( .A1(n11767), .A2(n18803), .B1(n11771), .Y(n18802) );
  xor2_1 U18447 ( .A(n18034), .B(n18804), .X(n11771) );
  nor2_1 U18448 ( .A(n11769), .B(n11770), .Y(n18804) );
  nand2_1 U18449 ( .A(n11769), .B(n11770), .Y(n18803) );
  xnor2_1 U18450 ( .A(n18805), .B(n18806), .Y(n11770) );
  xor2_1 U18451 ( .A(n18783), .B(n18792), .X(n18806) );
  xor2_1 U18452 ( .A(n24045), .B(n18807), .X(n18792) );
  a21oi_1 U18453 ( .A1(n11687), .A2(n18808), .B1(n18120), .Y(n18807) );
  nand2_1 U18454 ( .A(outData[30]), .B(n18124), .Y(n18808) );
  inv_1 U18455 ( .A(n11697), .Y(n18783) );
  xor2_1 U18456 ( .A(n18801), .B(n18809), .X(n11697) );
  xor2_1 U18457 ( .A(outData[31]), .B(n18800), .X(n18809) );
  inv_1 U18458 ( .A(n18798), .Y(n18800) );
  o22ai_1 U18459 ( .A1(n18810), .A2(n18811), .B1(n18124), .B2(n18812), .Y(
        n18798) );
  xor2_1 U18460 ( .A(n11677), .B(n18788), .X(n18805) );
  inv_1 U18461 ( .A(n18813), .Y(n18788) );
  o21ai_0 U18462 ( .A1(n18814), .A2(n18815), .B1(n18816), .Y(n18813) );
  xor2_1 U18463 ( .A(n18379), .B(n18817), .X(n18815) );
  xnor2_1 U18464 ( .A(n18818), .B(n18819), .Y(n11769) );
  xor2_1 U18465 ( .A(n17992), .B(n18820), .X(n18819) );
  xor2_1 U18466 ( .A(n11489), .B(n12476), .X(n18820) );
  xor2_1 U18467 ( .A(n11755), .B(n18821), .X(n18818) );
  xnor2_1 U18468 ( .A(n18822), .B(n12968), .Y(n11767) );
  a21oi_1 U18469 ( .A1(n11475), .A2(n11479), .B1(n11478), .Y(n18822) );
  xor2_1 U18470 ( .A(n12629), .B(n18823), .X(n11478) );
  nor2_1 U18471 ( .A(n18824), .B(n18825), .Y(n18823) );
  nand2_1 U18472 ( .A(n18824), .B(n18825), .Y(n11479) );
  xor2_1 U18473 ( .A(n18826), .B(n18827), .X(n18825) );
  nor2_1 U18474 ( .A(n18828), .B(n18829), .Y(n18827) );
  xor2_1 U18475 ( .A(n18814), .B(n18830), .X(n18824) );
  xor2_1 U18476 ( .A(n16742), .B(n18831), .X(n18830) );
  nand2_1 U18477 ( .A(n18816), .B(n18832), .Y(n18831) );
  inv_1 U18478 ( .A(n18817), .Y(n18832) );
  nor2_1 U18479 ( .A(n18833), .B(n18834), .Y(n18817) );
  nand2_1 U18480 ( .A(n18834), .B(n18833), .Y(n18816) );
  o22ai_1 U18481 ( .A1(n18835), .A2(n12958), .B1(n18836), .B2(n11746), .Y(
        n18833) );
  and2_0 U18482 ( .A(n18835), .B(n12958), .X(n18836) );
  inv_1 U18483 ( .A(n12953), .Y(n12958) );
  xor2_1 U18484 ( .A(n11687), .B(n18837), .X(n18834) );
  xnor2_1 U18485 ( .A(n18838), .B(n18839), .Y(n11687) );
  xor2_1 U18486 ( .A(n18812), .B(n18811), .X(n18839) );
  xor2_1 U18487 ( .A(n18840), .B(outData[31]), .X(n18838) );
  inv_1 U18488 ( .A(n17595), .Y(n16742) );
  nor4_1 U18489 ( .A(n18841), .B(n18842), .C(n18843), .D(n18844), .Y(n17595)
         );
  a21oi_1 U18490 ( .A1(n18845), .A2(n16188), .B1(n16171), .Y(n18842) );
  xor2_1 U18491 ( .A(n18846), .B(n17340), .X(n18814) );
  o22ai_1 U18492 ( .A1(n18847), .A2(n18848), .B1(n18849), .B2(n18850), .Y(
        n18846) );
  nor2_1 U18493 ( .A(n18851), .B(n18852), .Y(n18850) );
  inv_1 U18494 ( .A(n18851), .Y(n18848) );
  inv_1 U18495 ( .A(n18852), .Y(n18847) );
  o21ai_0 U18496 ( .A1(n18853), .A2(n11637), .B1(n11641), .Y(n11475) );
  xor2_1 U18497 ( .A(n10920), .B(n18854), .X(n11641) );
  and2_0 U18498 ( .A(n11640), .B(n11639), .X(n18854) );
  a21oi_1 U18499 ( .A1(n11651), .A2(n11652), .B1(n18855), .Y(n11637) );
  xnor2_1 U18500 ( .A(n18521), .B(n18856), .Y(n18855) );
  nand2_1 U18501 ( .A(n11646), .B(n18857), .Y(n18856) );
  inv_1 U18502 ( .A(n11653), .Y(n18857) );
  nor2_1 U18503 ( .A(n11651), .B(n11652), .Y(n11653) );
  o22ai_1 U18504 ( .A1(n12920), .A2(n12919), .B1(n18858), .B2(n12921), .Y(
        n11646) );
  o22ai_1 U18505 ( .A1(n11660), .A2(n11659), .B1(n18859), .B2(n11657), .Y(
        n12921) );
  xor2_1 U18506 ( .A(n18860), .B(n18861), .X(n11657) );
  nor2_1 U18507 ( .A(n18862), .B(n18863), .Y(n18861) );
  and2_0 U18508 ( .A(n11659), .B(n11660), .X(n18859) );
  xnor2_1 U18509 ( .A(n18864), .B(n12297), .Y(n11659) );
  o22ai_1 U18510 ( .A1(n18865), .A2(n18866), .B1(n18867), .B2(n11397), .Y(
        n18864) );
  xnor2_1 U18511 ( .A(n18868), .B(n18869), .Y(n11397) );
  xor2_1 U18512 ( .A(n18870), .B(n18111), .X(n18869) );
  xor2_1 U18513 ( .A(n11668), .B(n12515), .X(n18868) );
  nand4_1 U18514 ( .A(n18871), .B(n12409), .C(n18872), .D(n18873), .Y(n11668)
         );
  and2_0 U18515 ( .A(n12385), .B(n18874), .X(n18872) );
  nand3_1 U18516 ( .A(n24035), .B(n12383), .C(n24031), .Y(n18871) );
  nor2_1 U18517 ( .A(n11398), .B(n11399), .Y(n18867) );
  inv_1 U18518 ( .A(n18865), .Y(n11399) );
  inv_1 U18519 ( .A(n11398), .Y(n18866) );
  xor2_1 U18520 ( .A(n18875), .B(n18876), .X(n11398) );
  xor2_1 U18521 ( .A(n18040), .B(n18877), .X(n18876) );
  xnor2_1 U18522 ( .A(n18878), .B(n18879), .Y(n18875) );
  xor2_1 U18523 ( .A(n18880), .B(n17758), .X(n18865) );
  nand2_1 U18524 ( .A(n12561), .B(n12560), .Y(n18880) );
  nand2_1 U18525 ( .A(n12562), .B(n12557), .Y(n12560) );
  nand2_1 U18526 ( .A(n18881), .B(n18882), .Y(n12557) );
  inv_1 U18527 ( .A(n11429), .Y(n18882) );
  xnor2_1 U18528 ( .A(n18883), .B(n10919), .Y(n11429) );
  nand2_1 U18529 ( .A(n18884), .B(n18885), .Y(n18883) );
  xor2_1 U18530 ( .A(n18129), .B(n11430), .X(n18881) );
  nand2_1 U18531 ( .A(n11432), .B(n18886), .Y(n11430) );
  inv_1 U18532 ( .A(n11433), .Y(n18886) );
  nor2_1 U18533 ( .A(n18885), .B(n18884), .Y(n11433) );
  inv_1 U18534 ( .A(n18887), .Y(n18884) );
  o21ai_0 U18535 ( .A1(n1520), .A2(n18888), .B1(n18889), .Y(n18887) );
  mux2i_1 U18536 ( .A0(n18890), .A1(n18891), .S(n18892), .Y(n18889) );
  nor2_1 U18537 ( .A(n12901), .B(n10623), .Y(n18890) );
  xor2_1 U18538 ( .A(n18893), .B(n12901), .X(n18888) );
  inv_1 U18539 ( .A(n16637), .Y(n12901) );
  xnor2_1 U18540 ( .A(n18894), .B(n18895), .Y(n18885) );
  xnor2_1 U18541 ( .A(n18896), .B(n18897), .Y(n18895) );
  o22ai_1 U18542 ( .A1(n11448), .A2(n11449), .B1(n18898), .B2(n11446), .Y(
        n11432) );
  xnor2_1 U18543 ( .A(n18899), .B(n18900), .Y(n11446) );
  xor2_1 U18544 ( .A(n16823), .B(n18901), .X(n18900) );
  xor2_1 U18545 ( .A(n18902), .B(n18903), .X(n18899) );
  and2_0 U18546 ( .A(n11449), .B(n11448), .X(n18898) );
  xnor2_1 U18547 ( .A(n18904), .B(n18905), .Y(n11449) );
  nand2_1 U18548 ( .A(n18906), .B(n18907), .Y(n18904) );
  inv_1 U18549 ( .A(n18908), .Y(n18906) );
  nor2_1 U18550 ( .A(n11241), .B(n11246), .Y(n11448) );
  nor2_1 U18551 ( .A(n11245), .B(n18909), .Y(n11246) );
  inv_1 U18552 ( .A(n11244), .Y(n18909) );
  o21ai_0 U18553 ( .A1(n11254), .A2(n11255), .B1(n18910), .Y(n11244) );
  xor2_1 U18554 ( .A(n16246), .B(n18911), .X(n18910) );
  nand2_1 U18555 ( .A(n11252), .B(n11256), .Y(n18911) );
  nand2_1 U18556 ( .A(n11254), .B(n11255), .Y(n11256) );
  nand2_1 U18557 ( .A(n18912), .B(n11262), .Y(n11252) );
  nand2_1 U18558 ( .A(n18913), .B(n18914), .Y(n11262) );
  inv_1 U18559 ( .A(n18915), .Y(n18914) );
  xor2_1 U18560 ( .A(n18916), .B(n18917), .X(n18913) );
  xor2_1 U18561 ( .A(n17458), .B(n18918), .X(n18912) );
  nand2_1 U18562 ( .A(n11260), .B(n11261), .Y(n18918) );
  nand2_1 U18563 ( .A(n18915), .B(n18919), .Y(n11261) );
  xor2_1 U18564 ( .A(n18920), .B(n18916), .X(n18919) );
  nand2_1 U18565 ( .A(n18921), .B(n18922), .Y(n18916) );
  xor2_1 U18566 ( .A(n18923), .B(n18924), .X(n18915) );
  xor2_1 U18567 ( .A(n17766), .B(n18925), .X(n18924) );
  inv_1 U18568 ( .A(n16550), .Y(n17766) );
  xor2_1 U18569 ( .A(n11131), .B(n23676), .X(n18923) );
  inv_1 U18570 ( .A(n16757), .Y(n11131) );
  inv_1 U18571 ( .A(n18926), .Y(n11260) );
  o22ai_1 U18572 ( .A1(n11235), .A2(n11232), .B1(n18927), .B2(n11234), .Y(
        n18926) );
  o22ai_1 U18573 ( .A1(n11193), .A2(n11194), .B1(n18928), .B2(n18929), .Y(
        n11234) );
  and2_0 U18574 ( .A(n11194), .B(n11193), .X(n18929) );
  inv_1 U18575 ( .A(n11195), .Y(n18928) );
  o21ai_0 U18576 ( .A1(n18930), .A2(n11206), .B1(n11208), .Y(n11195) );
  nand2_1 U18577 ( .A(n18931), .B(n18932), .Y(n11208) );
  o22ai_1 U18578 ( .A1(n11282), .A2(n11285), .B1(n18933), .B2(n11283), .Y(
        n11206) );
  xnor2_1 U18579 ( .A(n18934), .B(n18935), .Y(n11283) );
  xnor2_1 U18580 ( .A(n18936), .B(n18937), .Y(n18935) );
  and2_0 U18581 ( .A(n11285), .B(n11282), .X(n18933) );
  xnor2_1 U18582 ( .A(n18938), .B(n13307), .Y(n11285) );
  o22ai_1 U18583 ( .A1(n18939), .A2(n11188), .B1(n18940), .B2(n11187), .Y(
        n18938) );
  xnor2_1 U18584 ( .A(n18941), .B(n18942), .Y(n11187) );
  xor2_1 U18585 ( .A(n18943), .B(n18944), .X(n18941) );
  and2_0 U18586 ( .A(n11188), .B(n18939), .X(n18940) );
  xnor2_1 U18587 ( .A(n18945), .B(n18946), .Y(n11188) );
  xor2_1 U18588 ( .A(n18947), .B(n18948), .X(n18946) );
  xor2_1 U18589 ( .A(n13368), .B(n23857), .X(n18948) );
  xor2_1 U18590 ( .A(n18949), .B(n11386), .X(n18945) );
  inv_1 U18591 ( .A(n16482), .Y(n11386) );
  inv_1 U18592 ( .A(n11186), .Y(n18939) );
  o22ai_1 U18593 ( .A1(n11144), .A2(n11146), .B1(n18950), .B2(n11145), .Y(
        n11186) );
  xor2_1 U18594 ( .A(n18951), .B(n12705), .X(n11145) );
  xor2_1 U18595 ( .A(n18952), .B(n23767), .X(n18951) );
  and2_0 U18596 ( .A(n11146), .B(n11144), .X(n18950) );
  xnor2_1 U18597 ( .A(n18953), .B(n18954), .Y(n11146) );
  xor2_1 U18598 ( .A(n18213), .B(n18955), .X(n18954) );
  xor2_1 U18599 ( .A(n18956), .B(n18957), .X(n18953) );
  xnor2_1 U18600 ( .A(n18958), .B(n18204), .Y(n11144) );
  nand2_1 U18601 ( .A(n18959), .B(n18960), .Y(n18958) );
  inv_1 U18602 ( .A(n11322), .Y(n18960) );
  xor2_1 U18603 ( .A(n12968), .B(n18961), .X(n11322) );
  nor2_1 U18604 ( .A(n11326), .B(n11327), .Y(n18961) );
  xor2_1 U18605 ( .A(n11328), .B(n18458), .X(n18959) );
  a21oi_1 U18606 ( .A1(n11327), .A2(n11326), .B1(n18962), .Y(n11328) );
  inv_1 U18607 ( .A(n11325), .Y(n18962) );
  xor2_1 U18608 ( .A(n16902), .B(n18963), .X(n11325) );
  a21oi_1 U18609 ( .A1(n12502), .A2(n12500), .B1(n18964), .Y(n18963) );
  inv_1 U18610 ( .A(n12503), .Y(n18964) );
  nand2_1 U18611 ( .A(n18965), .B(n18966), .Y(n12503) );
  o21ai_0 U18612 ( .A1(n11338), .A2(n11339), .B1(n18967), .Y(n12500) );
  xor2_1 U18613 ( .A(n18968), .B(n18969), .X(n18967) );
  nand2_1 U18614 ( .A(n11337), .B(n11340), .Y(n18969) );
  nand2_1 U18615 ( .A(n11338), .B(n11339), .Y(n11340) );
  o21ai_0 U18616 ( .A1(n12738), .A2(n12739), .B1(n18970), .Y(n11337) );
  xor2_1 U18617 ( .A(n17403), .B(n18971), .X(n18970) );
  nand2_1 U18618 ( .A(n12740), .B(n12736), .Y(n18971) );
  o22ai_1 U18619 ( .A1(n11540), .A2(n11541), .B1(n18972), .B2(n11538), .Y(
        n12736) );
  xnor2_1 U18620 ( .A(n18973), .B(n18974), .Y(n11538) );
  xor2_1 U18621 ( .A(n16940), .B(n18975), .X(n18974) );
  xor2_1 U18622 ( .A(n17598), .B(n23867), .X(n18973) );
  and2_0 U18623 ( .A(n11541), .B(n11540), .X(n18972) );
  xor2_1 U18624 ( .A(n18976), .B(n18977), .X(n11541) );
  xor2_1 U18625 ( .A(n18978), .B(n18979), .X(n18977) );
  a21oi_1 U18626 ( .A1(n17730), .A2(n18980), .B1(n18981), .Y(n11540) );
  inv_1 U18627 ( .A(n17729), .Y(n18981) );
  xor2_1 U18628 ( .A(n16750), .B(n18982), .X(n17729) );
  nor2_1 U18629 ( .A(n18983), .B(n18984), .Y(n18982) );
  inv_1 U18630 ( .A(n17726), .Y(n18980) );
  o22ai_1 U18631 ( .A1(n11562), .A2(n11564), .B1(n11565), .B2(n18985), .Y(
        n17726) );
  and2_0 U18632 ( .A(n11564), .B(n11562), .X(n18985) );
  inv_1 U18633 ( .A(n18986), .Y(n11565) );
  o21ai_0 U18634 ( .A1(n18987), .A2(n18988), .B1(n18989), .Y(n18986) );
  mux2i_1 U18635 ( .A0(n18990), .A1(n18991), .S(n18992), .Y(n18989) );
  nor2_1 U18636 ( .A(n18993), .B(n18994), .Y(n18991) );
  xor2_1 U18637 ( .A(n18992), .B(n18993), .X(n18988) );
  o22ai_1 U18638 ( .A1(n18995), .A2(n18996), .B1(n12799), .B2(n12795), .Y(
        n11564) );
  mux2i_1 U18639 ( .A0(n18997), .A1(n18998), .S(n18999), .Y(n12795) );
  o22ai_1 U18640 ( .A1(n19000), .A2(n17013), .B1(n19001), .B2(n19002), .Y(
        n18998) );
  nor2_1 U18641 ( .A(n19003), .B(n19004), .Y(n19001) );
  inv_1 U18642 ( .A(n19003), .Y(n17013) );
  nand2_1 U18643 ( .A(n19003), .B(n17014), .Y(n18997) );
  xnor2_1 U18644 ( .A(n19002), .B(n19004), .Y(n17014) );
  inv_1 U18645 ( .A(n19000), .Y(n19004) );
  xor2_1 U18646 ( .A(n16947), .B(n19005), .X(n19000) );
  xor2_1 U18647 ( .A(n23882), .B(n19006), .X(n19005) );
  xor2_1 U18648 ( .A(n19007), .B(n19008), .X(n19002) );
  xor2_1 U18649 ( .A(n19009), .B(n19010), .X(n19008) );
  xor2_1 U18650 ( .A(n19011), .B(n19012), .X(n19007) );
  xnor2_1 U18651 ( .A(n19013), .B(n11601), .Y(n19003) );
  nand2_1 U18652 ( .A(n19014), .B(n19015), .Y(n19013) );
  xor2_1 U18653 ( .A(n16843), .B(n19016), .X(n19015) );
  nand4_1 U18654 ( .A(n19017), .B(n19018), .C(n19019), .D(n19020), .Y(n19016)
         );
  xor2_1 U18655 ( .A(n19021), .B(n19022), .X(n19020) );
  nand2_1 U18656 ( .A(n19023), .B(n19024), .Y(n19022) );
  xor2_1 U18657 ( .A(n19025), .B(n19026), .X(n19019) );
  xor2_1 U18658 ( .A(n19027), .B(n19028), .X(n19026) );
  xor2_1 U18659 ( .A(n19029), .B(n19030), .X(n19018) );
  xor2_1 U18660 ( .A(n19031), .B(n19032), .X(n19017) );
  xor2_1 U18661 ( .A(n19033), .B(n12297), .X(n19031) );
  nand2_1 U18662 ( .A(n19034), .B(n19035), .Y(n19033) );
  xor2_1 U18663 ( .A(n19036), .B(n16737), .X(n19014) );
  nand3_1 U18664 ( .A(n19037), .B(n19038), .C(n19039), .Y(n19036) );
  xor2_1 U18665 ( .A(n19040), .B(n23903), .X(n19039) );
  inv_1 U18666 ( .A(n18605), .Y(n19038) );
  xor2_1 U18667 ( .A(n17525), .B(n19041), .X(n12799) );
  nor2_1 U18668 ( .A(n12797), .B(n12798), .Y(n19041) );
  inv_1 U18669 ( .A(n18995), .Y(n12798) );
  inv_1 U18670 ( .A(n12797), .Y(n18996) );
  xor2_1 U18671 ( .A(n19042), .B(n19043), .X(n12797) );
  xor2_1 U18672 ( .A(n17408), .B(n18358), .X(n19043) );
  inv_1 U18673 ( .A(n23863), .Y(n17408) );
  xor2_1 U18674 ( .A(n11120), .B(n19044), .X(n19042) );
  xor2_1 U18675 ( .A(n19045), .B(n19046), .X(n18995) );
  xor2_1 U18676 ( .A(n19047), .B(n17746), .X(n19046) );
  xor2_1 U18677 ( .A(n19048), .B(n19049), .X(n19045) );
  xnor2_1 U18678 ( .A(n16415), .B(n19050), .Y(n11562) );
  xor2_1 U18679 ( .A(n23869), .B(n19051), .X(n19050) );
  nand2_1 U18680 ( .A(n18983), .B(n18984), .Y(n17730) );
  xnor2_1 U18681 ( .A(n19052), .B(n19053), .Y(n18984) );
  xor2_1 U18682 ( .A(n19054), .B(n19055), .X(n19052) );
  mux2_1 U18683 ( .A0(n19056), .A1(n19057), .S(n2122), .X(n18983) );
  xor2_1 U18684 ( .A(n19058), .B(n17996), .X(n19057) );
  inv_1 U18685 ( .A(n19059), .Y(n17996) );
  xor2_1 U18686 ( .A(n19058), .B(n16674), .X(n19056) );
  xnor2_1 U18687 ( .A(n18521), .B(n19060), .Y(n12740) );
  and2_0 U18688 ( .A(n12739), .B(n12738), .X(n19060) );
  xnor2_1 U18689 ( .A(n19061), .B(n19062), .Y(n12739) );
  nand2_1 U18690 ( .A(n19063), .B(n19064), .Y(n19061) );
  inv_1 U18691 ( .A(n19065), .Y(n19064) );
  xor2_1 U18692 ( .A(n19066), .B(n19067), .X(n12738) );
  xnor2_1 U18693 ( .A(n19068), .B(n19069), .Y(n19066) );
  xor2_1 U18694 ( .A(n19070), .B(n17783), .X(n11339) );
  inv_1 U18695 ( .A(n12725), .Y(n17783) );
  nand2_1 U18696 ( .A(n19071), .B(n19072), .Y(n19070) );
  inv_1 U18697 ( .A(n19073), .Y(n19072) );
  xor2_1 U18698 ( .A(n19074), .B(n19075), .X(n11338) );
  xnor2_1 U18699 ( .A(n17152), .B(n19076), .Y(n19075) );
  xor2_1 U18700 ( .A(n19077), .B(n19078), .X(n19074) );
  xor2_1 U18701 ( .A(n11510), .B(n19079), .X(n12502) );
  nor2_1 U18702 ( .A(n18965), .B(n18966), .Y(n19079) );
  xnor2_1 U18703 ( .A(n19080), .B(n19081), .Y(n18966) );
  xor2_1 U18704 ( .A(n19082), .B(n23903), .X(n19080) );
  nand2_1 U18705 ( .A(n19083), .B(n19084), .Y(n19082) );
  xor2_1 U18706 ( .A(n19085), .B(n19086), .X(n18965) );
  xor2_1 U18707 ( .A(n23865), .B(n16933), .X(n19086) );
  inv_1 U18708 ( .A(n16707), .Y(n16902) );
  o221ai_1 U18709 ( .A1(n19087), .A2(n16187), .B1(n16141), .B2(n19088), .C1(
        n16184), .Y(n16707) );
  xor2_1 U18710 ( .A(n19089), .B(n19090), .X(n11326) );
  xor2_1 U18711 ( .A(n19091), .B(n19092), .X(n19089) );
  xnor2_1 U18712 ( .A(n19093), .B(n19094), .Y(n11327) );
  xor2_1 U18713 ( .A(n23864), .B(n18477), .X(n19094) );
  xor2_1 U18714 ( .A(n19095), .B(n12715), .X(n19093) );
  xnor2_1 U18715 ( .A(n19096), .B(n16507), .Y(n11282) );
  xor2_1 U18716 ( .A(n19097), .B(n12442), .X(n19096) );
  xor2_1 U18717 ( .A(n18125), .B(n11210), .X(n18930) );
  nor2_1 U18718 ( .A(n18931), .B(n18932), .Y(n11210) );
  xnor2_1 U18719 ( .A(n19098), .B(n19099), .Y(n18932) );
  xor2_1 U18720 ( .A(n19100), .B(n17697), .X(n19098) );
  nand2_1 U18721 ( .A(n19101), .B(n19102), .Y(n19100) );
  xor2_1 U18722 ( .A(n19103), .B(n16921), .X(n18931) );
  nand2_1 U18723 ( .A(n19104), .B(n19105), .Y(n19103) );
  inv_1 U18724 ( .A(n19106), .Y(n19104) );
  xor2_1 U18725 ( .A(n19107), .B(n19108), .X(n11194) );
  nand2_1 U18726 ( .A(n19109), .B(n19110), .Y(n19107) );
  inv_1 U18727 ( .A(n19111), .Y(n19109) );
  xor2_1 U18728 ( .A(n19112), .B(n19113), .X(n11193) );
  xor2_1 U18729 ( .A(n19114), .B(n19115), .X(n19112) );
  and2_0 U18730 ( .A(n11232), .B(n11235), .X(n18927) );
  xnor2_1 U18731 ( .A(n19116), .B(n19117), .Y(n11232) );
  xnor2_1 U18732 ( .A(n19118), .B(n19119), .Y(n19116) );
  nor2_1 U18733 ( .A(n19120), .B(n19121), .Y(n11235) );
  a21oi_1 U18734 ( .A1(n19122), .A2(n19123), .B1(n19124), .Y(n19120) );
  xnor2_1 U18735 ( .A(n19125), .B(n19126), .Y(n11255) );
  xor2_1 U18736 ( .A(n2116), .B(n11751), .X(n19126) );
  xor2_1 U18737 ( .A(n19127), .B(n16906), .X(n19125) );
  xor2_1 U18738 ( .A(n19128), .B(n19129), .X(n11254) );
  xnor2_1 U18739 ( .A(n19130), .B(n19131), .Y(n19129) );
  xor2_1 U18740 ( .A(n19132), .B(n11520), .X(n19128) );
  xor2_1 U18741 ( .A(n19133), .B(n16829), .X(n11245) );
  nand2_1 U18742 ( .A(n19134), .B(n19135), .Y(n19133) );
  nor2_1 U18743 ( .A(n19135), .B(n19134), .Y(n11241) );
  xnor2_1 U18744 ( .A(n19136), .B(n19137), .Y(n19134) );
  xor2_1 U18745 ( .A(n19138), .B(n19139), .X(n19136) );
  xor2_1 U18746 ( .A(n19140), .B(n19141), .X(n19135) );
  xor2_1 U18747 ( .A(n23702), .B(n16737), .X(n19141) );
  nor4_1 U18748 ( .A(n19142), .B(n19143), .C(n19144), .D(n19145), .Y(n16737)
         );
  o32ai_1 U18749 ( .A1(n14696), .A2(n24046), .A3(n24038), .B1(n14665), .B2(
        n14663), .Y(n19145) );
  a21oi_1 U18750 ( .A1(n14625), .A2(n14694), .B1(n24039), .Y(n19144) );
  nand2_1 U18751 ( .A(n19146), .B(n14676), .Y(n14694) );
  a21oi_1 U18752 ( .A1(n14699), .A2(n14695), .B1(n14707), .Y(n19143) );
  xor2_1 U18753 ( .A(n19147), .B(n17761), .X(n19140) );
  inv_1 U18754 ( .A(n12942), .Y(n18129) );
  nand2_1 U18755 ( .A(n19148), .B(n19149), .Y(n12562) );
  xor2_1 U18756 ( .A(n17765), .B(n19150), .X(n19148) );
  nand2_1 U18757 ( .A(n19151), .B(n19150), .Y(n12561) );
  inv_1 U18758 ( .A(n19152), .Y(n19150) );
  o21ai_0 U18759 ( .A1(n12894), .A2(n19153), .B1(n19154), .Y(n19152) );
  mux2i_1 U18760 ( .A0(n19155), .A1(n19156), .S(n19157), .Y(n19154) );
  nor2_1 U18761 ( .A(n8), .B(n12890), .Y(n19155) );
  xor2_1 U18762 ( .A(n19157), .B(n16894), .X(n19153) );
  xor2_1 U18763 ( .A(n12297), .B(n19149), .X(n19151) );
  o21ai_0 U18764 ( .A1(n19158), .A2(n19159), .B1(n19160), .Y(n19149) );
  mux2i_1 U18765 ( .A0(n19161), .A1(n19162), .S(n19163), .Y(n19160) );
  nor2_1 U18766 ( .A(n19164), .B(n19165), .Y(n19162) );
  xor2_1 U18767 ( .A(n19163), .B(n19165), .X(n19159) );
  xnor2_1 U18768 ( .A(n19166), .B(n19167), .Y(n19163) );
  xor2_1 U18769 ( .A(n16535), .B(n19168), .X(n19167) );
  xor2_1 U18770 ( .A(n19169), .B(n19170), .X(n11660) );
  xor2_1 U18771 ( .A(n17003), .B(n1519), .X(n19169) );
  and2_0 U18772 ( .A(n12919), .B(n12920), .X(n18858) );
  xor2_1 U18773 ( .A(n19171), .B(n19172), .X(n12919) );
  xor2_1 U18774 ( .A(n19173), .B(n19174), .X(n19172) );
  xnor2_1 U18775 ( .A(n19175), .B(n19176), .Y(n12920) );
  xor2_1 U18776 ( .A(n12445), .B(n12297), .X(n19176) );
  nand2_1 U18777 ( .A(n19177), .B(n19178), .Y(n19175) );
  inv_1 U18778 ( .A(n19179), .Y(n19178) );
  xnor2_1 U18779 ( .A(n19180), .B(n16307), .Y(n11652) );
  xor2_1 U18780 ( .A(n12446), .B(n19181), .X(n19180) );
  xnor2_1 U18781 ( .A(n19182), .B(n19183), .Y(n11651) );
  xor2_1 U18782 ( .A(n17992), .B(n19184), .X(n19183) );
  nand2_1 U18783 ( .A(n19185), .B(n19186), .Y(n19184) );
  inv_1 U18784 ( .A(n19187), .Y(n19185) );
  nor2_1 U18785 ( .A(n11639), .B(n11640), .Y(n18853) );
  xnor2_1 U18786 ( .A(n19188), .B(n19189), .Y(n11640) );
  xor2_1 U18787 ( .A(n18851), .B(n18852), .X(n19189) );
  mux2i_1 U18788 ( .A0(n19190), .A1(n19191), .S(n17746), .Y(n18852) );
  mux2i_1 U18789 ( .A0(n19192), .A1(n19193), .S(n18476), .Y(n19191) );
  nand2_1 U18790 ( .A(n19194), .B(n19195), .Y(n19193) );
  o22ai_1 U18791 ( .A1(n19196), .A2(n18476), .B1(n19197), .B2(n19194), .Y(
        n19190) );
  inv_1 U18792 ( .A(n19192), .Y(n19196) );
  xor2_1 U18793 ( .A(n19198), .B(n19199), .X(n18851) );
  xor2_1 U18794 ( .A(n11746), .B(n19200), .X(n19199) );
  inv_1 U18795 ( .A(n11570), .Y(n19200) );
  xor2_1 U18796 ( .A(n18835), .B(n12953), .X(n19198) );
  o22ai_1 U18797 ( .A1(n19201), .A2(n18812), .B1(outData[31]), .B2(n19202), 
        .Y(n12953) );
  a21oi_1 U18798 ( .A1(n19203), .A2(n19204), .B1(n19205), .Y(n19202) );
  o21ai_0 U18799 ( .A1(n19206), .A2(n19207), .B1(n19205), .Y(n18812) );
  inv_1 U18800 ( .A(n18810), .Y(n19205) );
  nor2_1 U18801 ( .A(n19201), .B(outData[31]), .Y(n18810) );
  inv_1 U18802 ( .A(n19204), .Y(n19206) );
  nor2_1 U18803 ( .A(n19204), .B(n19203), .Y(n19201) );
  inv_1 U18804 ( .A(n19207), .Y(n19203) );
  o21ai_0 U18805 ( .A1(n10930), .A2(n19208), .B1(n19209), .Y(n19204) );
  xor2_1 U18806 ( .A(n12297), .B(n19210), .X(n19209) );
  nor2_1 U18807 ( .A(n19211), .B(n19212), .Y(n19210) );
  xor2_1 U18808 ( .A(n12821), .B(n18849), .X(n19188) );
  inv_1 U18809 ( .A(n19213), .Y(n18849) );
  o21ai_0 U18810 ( .A1(n19182), .A2(n19214), .B1(n19186), .Y(n19213) );
  nand2_1 U18811 ( .A(n19215), .B(n19216), .Y(n19186) );
  xor2_1 U18812 ( .A(n11684), .B(n19187), .X(n19214) );
  nor2_1 U18813 ( .A(n19216), .B(n19215), .Y(n19187) );
  xnor2_1 U18814 ( .A(n19217), .B(n18476), .Y(n19215) );
  inv_1 U18815 ( .A(n18473), .Y(n18476) );
  o21ai_0 U18816 ( .A1(n19208), .A2(n19218), .B1(n19219), .Y(n18473) );
  mux2i_1 U18817 ( .A0(n19220), .A1(n19211), .S(n19212), .Y(n19219) );
  inv_1 U18818 ( .A(n19221), .Y(n19212) );
  and2_0 U18819 ( .A(n10930), .B(n19208), .X(n19211) );
  nor2_1 U18820 ( .A(n19222), .B(n10930), .Y(n19220) );
  xor2_1 U18821 ( .A(n19221), .B(n10930), .X(n19218) );
  xnor2_1 U18822 ( .A(n18837), .B(n19223), .Y(n10930) );
  a21oi_1 U18823 ( .A1(n19224), .A2(n19225), .B1(n18835), .Y(n19223) );
  nor2_1 U18824 ( .A(n11498), .B(outData[31]), .Y(n18835) );
  nand2_1 U18825 ( .A(outData[31]), .B(n11498), .Y(n19225) );
  a21oi_1 U18826 ( .A1(n18124), .A2(outData[30]), .B1(n18120), .Y(n18837) );
  nor2_1 U18827 ( .A(n18124), .B(outData[30]), .Y(n18120) );
  inv_1 U18828 ( .A(outData[31]), .Y(n18124) );
  o21ai_0 U18829 ( .A1(n19226), .A2(n18779), .B1(n19227), .Y(n19221) );
  xor2_1 U18830 ( .A(n13009), .B(n19228), .X(n19227) );
  nor2_1 U18831 ( .A(n19229), .B(n19230), .Y(n19228) );
  o21ai_0 U18832 ( .A1(n19197), .A2(n19194), .B1(n19192), .Y(n19217) );
  nand2_1 U18833 ( .A(n19197), .B(n19194), .Y(n19192) );
  inv_1 U18834 ( .A(n19195), .Y(n19197) );
  o21ai_0 U18835 ( .A1(n19231), .A2(n11681), .B1(n19232), .Y(n19216) );
  xnor2_1 U18836 ( .A(n11601), .B(n19233), .Y(n19232) );
  o221ai_1 U18837 ( .A1(n19234), .A2(n13950), .B1(n19235), .B2(n19236), .C1(
        n19237), .Y(n11601) );
  nor2_1 U18838 ( .A(n19238), .B(n19239), .Y(n19237) );
  xor2_1 U18839 ( .A(n19240), .B(n19241), .X(n19182) );
  o21ai_0 U18840 ( .A1(n19242), .A2(n19243), .B1(n19244), .Y(n19240) );
  xnor2_1 U18841 ( .A(n19245), .B(n16843), .Y(n19244) );
  nand2_1 U18842 ( .A(n19171), .B(n19173), .Y(n19245) );
  inv_1 U18843 ( .A(n19174), .Y(n19243) );
  o21ai_0 U18844 ( .A1(n18860), .A2(n19246), .B1(n19247), .Y(n19174) );
  xor2_1 U18845 ( .A(n10942), .B(n18862), .X(n19247) );
  and2_0 U18846 ( .A(n19248), .B(n19249), .X(n18862) );
  xor2_1 U18847 ( .A(n11520), .B(n18863), .X(n19246) );
  nor2_1 U18848 ( .A(n19249), .B(n19248), .Y(n18863) );
  xnor2_1 U18849 ( .A(n18486), .B(n19250), .Y(n19248) );
  a21oi_1 U18850 ( .A1(n19251), .A2(n19252), .B1(n19253), .Y(n19250) );
  inv_1 U18851 ( .A(n12938), .Y(n18486) );
  nand2_1 U18852 ( .A(n19254), .B(n19255), .Y(n19249) );
  o21ai_0 U18853 ( .A1(n19256), .A2(n19257), .B1(n19258), .Y(n19255) );
  inv_1 U18854 ( .A(n19259), .Y(n19256) );
  xor2_1 U18855 ( .A(n18532), .B(n19260), .X(n19254) );
  nor2_1 U18856 ( .A(n19259), .B(n18491), .Y(n19260) );
  inv_1 U18857 ( .A(n19257), .Y(n18491) );
  a21oi_1 U18858 ( .A1(n18877), .A2(n18879), .B1(n19261), .Y(n18860) );
  xor2_1 U18859 ( .A(n18968), .B(n19262), .X(n19261) );
  nor2_1 U18860 ( .A(n19263), .B(n18878), .Y(n19262) );
  xnor2_1 U18861 ( .A(n13401), .B(n19264), .Y(n18878) );
  a21oi_1 U18862 ( .A1(n19265), .A2(n19166), .B1(n19161), .Y(n19264) );
  nor2_1 U18863 ( .A(n19164), .B(n19266), .Y(n19161) );
  inv_1 U18864 ( .A(n19158), .Y(n19164) );
  o22ai_1 U18865 ( .A1(n18896), .A2(n18897), .B1(n19267), .B2(n18894), .Y(
        n19166) );
  xnor2_1 U18866 ( .A(n19268), .B(n12944), .Y(n18894) );
  xor2_1 U18867 ( .A(n19269), .B(n17915), .X(n19268) );
  nand2_1 U18868 ( .A(n19270), .B(n19271), .Y(n19269) );
  inv_1 U18869 ( .A(n19272), .Y(n19271) );
  and2_0 U18870 ( .A(n18897), .B(n18896), .X(n19267) );
  o22ai_1 U18871 ( .A1(n19273), .A2(n19274), .B1(n19275), .B2(n19276), .Y(
        n18897) );
  inv_1 U18872 ( .A(n19277), .Y(n19276) );
  nor2_1 U18873 ( .A(outData[24]), .B(outData[22]), .Y(n19275) );
  inv_1 U18874 ( .A(n17047), .Y(n19274) );
  a22oi_1 U18875 ( .A1(n18903), .A2(n18901), .B1(n18902), .B2(n19278), .Y(
        n18896) );
  xor2_1 U18876 ( .A(n18624), .B(n19279), .X(n19278) );
  nor2_1 U18877 ( .A(n18901), .B(n18903), .Y(n19279) );
  inv_1 U18878 ( .A(n17403), .Y(n18624) );
  o22ai_1 U18879 ( .A1(n19137), .A2(n19138), .B1(n19139), .B2(n19280), .Y(
        n18902) );
  and2_0 U18880 ( .A(n19138), .B(n19137), .X(n19280) );
  inv_1 U18881 ( .A(n19281), .Y(n19139) );
  o22ai_1 U18882 ( .A1(n11223), .A2(n19282), .B1(n19283), .B2(n19284), .Y(
        n19281) );
  and2_0 U18883 ( .A(n19282), .B(n11223), .X(n19283) );
  xor2_1 U18884 ( .A(n18505), .B(n19285), .X(n19138) );
  nor2_1 U18885 ( .A(n19286), .B(n19287), .Y(n19285) );
  inv_1 U18886 ( .A(n19288), .Y(n19286) );
  xor2_1 U18887 ( .A(n19289), .B(n18118), .X(n19137) );
  o21ai_0 U18888 ( .A1(n19131), .A2(n19130), .B1(n19290), .Y(n19289) );
  xor2_1 U18889 ( .A(n17506), .B(n19291), .X(n19290) );
  a21oi_1 U18890 ( .A1(n19131), .A2(n19130), .B1(n19132), .Y(n19291) );
  a21oi_1 U18891 ( .A1(n18921), .A2(n18917), .B1(n19292), .Y(n19132) );
  inv_1 U18892 ( .A(n18922), .Y(n19292) );
  nand2_1 U18893 ( .A(n19293), .B(n19294), .Y(n18922) );
  inv_1 U18894 ( .A(n18920), .Y(n18917) );
  o22ai_1 U18895 ( .A1(n18131), .A2(n18652), .B1(n19295), .B2(n12978), .Y(
        n18920) );
  and2_0 U18896 ( .A(n18131), .B(n18652), .X(n19295) );
  or2_0 U18897 ( .A(n19294), .B(n19293), .X(n18921) );
  xnor2_1 U18898 ( .A(n19296), .B(n19297), .Y(n19293) );
  xor2_1 U18899 ( .A(n18508), .B(n19298), .X(n19296) );
  o22ai_1 U18900 ( .A1(n19119), .A2(n19118), .B1(n19299), .B2(n19117), .Y(
        n19294) );
  xor2_1 U18901 ( .A(n19300), .B(n18652), .X(n19117) );
  xor2_1 U18902 ( .A(n19301), .B(n19302), .X(n18652) );
  xor2_1 U18903 ( .A(n11413), .B(n16535), .X(n19302) );
  xnor2_1 U18904 ( .A(n19303), .B(n19304), .Y(n19301) );
  nand2_1 U18905 ( .A(n19305), .B(n19306), .Y(n19303) );
  xnor2_1 U18906 ( .A(n18131), .B(n12978), .Y(n19300) );
  nor2_1 U18907 ( .A(outData[18]), .B(outData[20]), .Y(n18131) );
  and2_0 U18908 ( .A(n19118), .B(n19119), .X(n19299) );
  o22ai_1 U18909 ( .A1(n19307), .A2(n19308), .B1(n19309), .B2(n19113), .Y(
        n19118) );
  xnor2_1 U18910 ( .A(n19310), .B(n19311), .Y(n19113) );
  xnor2_1 U18911 ( .A(n19312), .B(n10796), .Y(n19311) );
  nand4_1 U18912 ( .A(n19313), .B(n19314), .C(n19315), .D(n12416), .Y(n10796)
         );
  nand2_1 U18913 ( .A(n19316), .B(n24030), .Y(n19314) );
  mux2_1 U18914 ( .A0(n19317), .A1(n19318), .S(n10610), .X(n19316) );
  mux2i_1 U18915 ( .A0(n19319), .A1(n12419), .S(n24027), .Y(n19313) );
  nor2_1 U18916 ( .A(n12370), .B(n10610), .Y(n19319) );
  xor2_1 U18917 ( .A(n18525), .B(n19320), .X(n19310) );
  nor2_1 U18918 ( .A(n19115), .B(n19114), .Y(n19309) );
  inv_1 U18919 ( .A(n19308), .Y(n19115) );
  o22ai_1 U18920 ( .A1(n11166), .A2(n19321), .B1(n19322), .B2(n19323), .Y(
        n19308) );
  inv_1 U18921 ( .A(n19324), .Y(n19323) );
  and2_0 U18922 ( .A(n19321), .B(n11166), .X(n19322) );
  inv_1 U18923 ( .A(n11163), .Y(n11166) );
  inv_1 U18924 ( .A(n19114), .Y(n19307) );
  xor2_1 U18925 ( .A(n11520), .B(n19325), .X(n19114) );
  a21oi_1 U18926 ( .A1(n19099), .A2(n19102), .B1(n19326), .Y(n19325) );
  xor2_1 U18927 ( .A(n19327), .B(n19101), .X(n19326) );
  nand2_1 U18928 ( .A(n19328), .B(n19329), .Y(n19101) );
  inv_1 U18929 ( .A(n19330), .Y(n19329) );
  xor2_1 U18930 ( .A(n17310), .B(n19331), .X(n19328) );
  nand2_1 U18931 ( .A(n19330), .B(n19332), .Y(n19102) );
  xor2_1 U18932 ( .A(n19331), .B(n12629), .X(n19332) );
  o22ai_1 U18933 ( .A1(n19333), .A2(n19334), .B1(n18537), .B2(n19335), .Y(
        n19331) );
  nor2_1 U18934 ( .A(n19336), .B(n19337), .Y(n19335) );
  xor2_1 U18935 ( .A(n18068), .B(n19334), .X(n19337) );
  a21oi_1 U18936 ( .A1(n18537), .A2(n19338), .B1(n19336), .Y(n19333) );
  inv_1 U18937 ( .A(n18642), .Y(n18537) );
  xor2_1 U18938 ( .A(n11163), .B(n19339), .X(n19330) );
  xor2_1 U18939 ( .A(n19324), .B(n19321), .X(n19339) );
  xnor2_1 U18940 ( .A(n17620), .B(n19340), .Y(n19321) );
  nor2_1 U18941 ( .A(outData[18]), .B(outData[16]), .Y(n19340) );
  mux2i_1 U18942 ( .A0(n19341), .A1(n19342), .S(n19343), .Y(n11163) );
  xor2_1 U18943 ( .A(n19344), .B(n19345), .X(n19342) );
  xor2_1 U18944 ( .A(n19344), .B(n19346), .X(n19341) );
  o22ai_1 U18945 ( .A1(n18934), .A2(n18937), .B1(n18936), .B2(n19347), .Y(
        n19099) );
  and2_0 U18946 ( .A(n18937), .B(n18934), .X(n19347) );
  and2_0 U18947 ( .A(n19348), .B(n19349), .X(n18936) );
  o21ai_0 U18948 ( .A1(n18944), .A2(n18943), .B1(n18942), .Y(n19349) );
  xnor2_1 U18949 ( .A(n19350), .B(n14685), .Y(n18942) );
  o22ai_1 U18950 ( .A1(n18957), .A2(n19351), .B1(n19352), .B2(n19353), .Y(
        n19350) );
  nor2_1 U18951 ( .A(n18956), .B(n19354), .Y(n19353) );
  inv_1 U18952 ( .A(n18955), .Y(n19352) );
  o22ai_1 U18953 ( .A1(n19090), .A2(n19355), .B1(n19356), .B2(n19357), .Y(
        n18955) );
  and2_0 U18954 ( .A(n19355), .B(n19090), .X(n19357) );
  inv_1 U18955 ( .A(n19091), .Y(n19356) );
  o22ai_1 U18956 ( .A1(n19358), .A2(n19359), .B1(n19360), .B2(n19361), .Y(
        n19091) );
  mux2i_1 U18957 ( .A0(n19362), .A1(n19363), .S(n18128), .Y(n19361) );
  nor2_1 U18958 ( .A(n19363), .B(n18555), .Y(n19362) );
  xor2_1 U18959 ( .A(n16763), .B(n19364), .X(n19359) );
  inv_1 U18960 ( .A(n19092), .Y(n19355) );
  a21oi_1 U18961 ( .A1(n19084), .A2(n19081), .B1(n19365), .Y(n19092) );
  inv_1 U18962 ( .A(n19083), .Y(n19365) );
  nand2_1 U18963 ( .A(n19366), .B(n19367), .Y(n19083) );
  xor2_1 U18964 ( .A(n19368), .B(n11414), .X(n19081) );
  o22ai_1 U18965 ( .A1(n19369), .A2(n19370), .B1(n19076), .B2(n19371), .Y(
        n19368) );
  nor2_1 U18966 ( .A(n19078), .B(n19077), .Y(n19371) );
  inv_1 U18967 ( .A(n19370), .Y(n19078) );
  nor2_1 U18968 ( .A(n19372), .B(n19373), .Y(n19076) );
  a21oi_1 U18969 ( .A1(n19068), .A2(n19067), .B1(n19069), .Y(n19373) );
  a21oi_1 U18970 ( .A1(n18978), .A2(n18976), .B1(n19374), .Y(n19069) );
  xor2_1 U18971 ( .A(n19375), .B(n19376), .X(n19374) );
  nand2_1 U18972 ( .A(n19377), .B(n18979), .Y(n19376) );
  o22ai_1 U18973 ( .A1(n19053), .A2(n19055), .B1(n19054), .B2(n19378), .Y(
        n18979) );
  and2_0 U18974 ( .A(n19055), .B(n19053), .X(n19378) );
  inv_1 U18975 ( .A(n19379), .Y(n19054) );
  o22ai_1 U18976 ( .A1(n18987), .A2(n18993), .B1(n18992), .B2(n19380), .Y(
        n19379) );
  xor2_1 U18977 ( .A(n17746), .B(n18990), .X(n19380) );
  and2_0 U18978 ( .A(n18987), .B(n18993), .X(n18990) );
  xor2_1 U18979 ( .A(n19381), .B(n19382), .X(n18992) );
  o22ai_1 U18980 ( .A1(n19383), .A2(n19047), .B1(n19384), .B2(n19048), .Y(
        n19381) );
  xnor2_1 U18981 ( .A(n19385), .B(n18588), .Y(n19048) );
  xor2_1 U18982 ( .A(n19386), .B(n19387), .X(n19385) );
  and2_0 U18983 ( .A(n19047), .B(n19383), .X(n19384) );
  o21ai_0 U18984 ( .A1(n19388), .A2(n19389), .B1(n19390), .Y(n19047) );
  inv_1 U18985 ( .A(n19049), .Y(n19383) );
  o22ai_1 U18986 ( .A1(n19391), .A2(n19011), .B1(n19392), .B2(n19012), .Y(
        n19049) );
  mux2i_1 U18987 ( .A0(n19393), .A1(n19394), .S(n11414), .Y(n19012) );
  o211ai_1 U18988 ( .A1(n10621), .A2(n19395), .B1(n13960), .C1(n19396), .Y(
        n11414) );
  nand2_1 U18989 ( .A(n19030), .B(n19397), .Y(n19394) );
  xor2_1 U18990 ( .A(n19398), .B(n19399), .X(n19030) );
  o22ai_1 U18991 ( .A1(n19029), .A2(n19398), .B1(n19400), .B2(n19399), .Y(
        n19393) );
  xor2_1 U18992 ( .A(n16757), .B(n19401), .X(n19399) );
  a222oi_1 U18993 ( .A1(n18611), .A2(n19402), .B1(n19403), .B2(n12968), .C1(
        n19404), .C2(n19405), .Y(n19401) );
  inv_1 U18994 ( .A(n19406), .Y(n19402) );
  a21oi_1 U18995 ( .A1(n19405), .A2(n23903), .B1(n19404), .Y(n19406) );
  a211oi_1 U18996 ( .A1(n19407), .A2(n19408), .B1(n18841), .C1(n19409), .Y(
        n16757) );
  inv_1 U18997 ( .A(n19410), .Y(n19409) );
  a222oi_1 U18998 ( .A1(n16107), .A2(n19411), .B1(n16124), .B2(n19412), .C1(
        n23975), .C2(n19413), .Y(n19410) );
  o22ai_1 U18999 ( .A1(n19407), .A2(n19414), .B1(n16171), .B2(n19415), .Y(
        n19413) );
  inv_1 U19000 ( .A(n16134), .Y(n16171) );
  nand2_1 U19001 ( .A(n18845), .B(n16121), .Y(n19412) );
  o21ai_0 U19002 ( .A1(n23978), .A2(n16139), .B1(n16178), .Y(n18841) );
  and2_0 U19003 ( .A(n19398), .B(n19029), .X(n19400) );
  xor2_1 U19004 ( .A(n19416), .B(n19417), .X(n19398) );
  nand2_1 U19005 ( .A(n19418), .B(n19419), .Y(n19416) );
  inv_1 U19006 ( .A(n19397), .Y(n19029) );
  o22ai_1 U19007 ( .A1(n19420), .A2(n19421), .B1(n19028), .B2(n19422), .Y(
        n19397) );
  nor2_1 U19008 ( .A(n19027), .B(n19025), .Y(n19422) );
  a21oi_1 U19009 ( .A1(n19021), .A2(n19423), .B1(n19424), .Y(n19028) );
  inv_1 U19010 ( .A(n19024), .Y(n19424) );
  nand2_1 U19011 ( .A(n19425), .B(n19426), .Y(n19024) );
  xor2_1 U19012 ( .A(n19023), .B(n18050), .X(n19423) );
  nand2_1 U19013 ( .A(n19427), .B(n16167), .Y(n18050) );
  o21ai_0 U19014 ( .A1(n16100), .A2(n16155), .B1(n19428), .Y(n19427) );
  nand4_1 U19015 ( .A(n19429), .B(n16166), .C(n16186), .D(n14215), .Y(n19428)
         );
  o21ai_0 U19016 ( .A1(n23962), .A2(n16168), .B1(n23964), .Y(n19429) );
  or2_0 U19017 ( .A(n19426), .B(n19425), .X(n19023) );
  inv_1 U19018 ( .A(n19430), .Y(n19425) );
  o21ai_0 U19019 ( .A1(n18607), .A2(n19431), .B1(n19432), .Y(n19430) );
  mux2i_1 U19020 ( .A0(n19433), .A1(n19434), .S(n19435), .Y(n19432) );
  nor2_1 U19021 ( .A(n19436), .B(n19437), .Y(n19433) );
  xor2_1 U19022 ( .A(n19435), .B(n19438), .X(n19431) );
  xor2_1 U19023 ( .A(n16773), .B(n19439), .X(n19435) );
  inv_1 U19024 ( .A(n18947), .Y(n16773) );
  o22ai_1 U19025 ( .A1(n19440), .A2(n18609), .B1(outData[2]), .B2(n19441), .Y(
        n19426) );
  nor2_1 U19026 ( .A(n19442), .B(n19443), .Y(n19441) );
  o21ai_0 U19027 ( .A1(n19444), .A2(n19032), .B1(n19035), .Y(n19021) );
  o211ai_1 U19028 ( .A1(n19445), .A2(n18606), .B1(n19446), .C1(n19447), .Y(
        n19035) );
  xnor2_1 U19029 ( .A(n18651), .B(n19448), .Y(n19032) );
  o21ai_0 U19030 ( .A1(n18605), .A2(n18138), .B1(n19037), .Y(n19448) );
  xor2_1 U19031 ( .A(n18606), .B(n19449), .X(n19037) );
  xor2_1 U19032 ( .A(n19168), .B(n19450), .X(n18605) );
  a21oi_1 U19033 ( .A1(n19449), .A2(n19040), .B1(n19451), .Y(n19450) );
  inv_1 U19034 ( .A(n19452), .Y(n19451) );
  xor2_1 U19035 ( .A(n19034), .B(n19453), .X(n19444) );
  inv_1 U19036 ( .A(n19454), .Y(n19034) );
  a211oi_1 U19037 ( .A1(n19446), .A2(n18606), .B1(n19445), .C1(n19447), .Y(
        n19454) );
  xnor2_1 U19038 ( .A(n19455), .B(n19443), .Y(n19447) );
  xor2_1 U19039 ( .A(n18609), .B(n12308), .X(n19455) );
  inv_1 U19040 ( .A(n19442), .Y(n18609) );
  a21oi_1 U19041 ( .A1(n19456), .A2(n19457), .B1(n19458), .Y(n19442) );
  and2_0 U19042 ( .A(n19459), .B(n19456), .X(n18606) );
  xor2_1 U19043 ( .A(n10893), .B(n19460), .X(n19459) );
  nand2_1 U19044 ( .A(n19452), .B(n19461), .Y(n19460) );
  inv_1 U19045 ( .A(n19027), .Y(n19421) );
  xnor2_1 U19046 ( .A(n19403), .B(n19404), .Y(n19027) );
  xor2_1 U19047 ( .A(n19462), .B(n17774), .X(n19404) );
  xor2_1 U19048 ( .A(n18611), .B(n19405), .X(n19403) );
  xor2_1 U19049 ( .A(n11103), .B(n19463), .X(n19405) );
  nor2_1 U19050 ( .A(outData[4]), .B(outData[2]), .Y(n19463) );
  xnor2_1 U19051 ( .A(n19464), .B(n19465), .Y(n18611) );
  xor2_1 U19052 ( .A(outData[0]), .B(n19466), .X(n19465) );
  xor2_1 U19053 ( .A(n19467), .B(n19468), .X(n19464) );
  inv_1 U19054 ( .A(n19025), .Y(n19420) );
  mux2i_1 U19055 ( .A0(n19469), .A1(n19470), .S(n17479), .Y(n19025) );
  o22ai_1 U19056 ( .A1(n19437), .A2(n18607), .B1(n19439), .B2(n19434), .Y(
        n19470) );
  inv_1 U19057 ( .A(n19471), .Y(n19434) );
  mux2i_1 U19058 ( .A0(n19471), .A1(n19472), .S(n19439), .Y(n19469) );
  nand2_1 U19059 ( .A(n19436), .B(n19437), .Y(n19472) );
  inv_1 U19060 ( .A(n18607), .Y(n19436) );
  nand2_1 U19061 ( .A(n19437), .B(n18607), .Y(n19471) );
  xor2_1 U19062 ( .A(n19473), .B(n16898), .X(n18607) );
  inv_1 U19063 ( .A(n10808), .Y(n16898) );
  nand4_1 U19064 ( .A(n19474), .B(n13898), .C(n13934), .D(n16148), .Y(n10808)
         );
  nand2_1 U19065 ( .A(n13926), .B(n13922), .Y(n13898) );
  nand2_1 U19066 ( .A(n13915), .B(n24000), .Y(n19474) );
  nand2_1 U19067 ( .A(n19475), .B(n19467), .Y(n19473) );
  xor2_1 U19068 ( .A(n12512), .B(n19476), .X(n19475) );
  nor2_1 U19069 ( .A(n19458), .B(n19477), .Y(n19476) );
  inv_1 U19070 ( .A(n19438), .Y(n19437) );
  xnor2_1 U19071 ( .A(outData[2]), .B(outData[4]), .Y(n19438) );
  and2_0 U19072 ( .A(n19011), .B(n19391), .X(n19392) );
  xor2_1 U19073 ( .A(n19478), .B(n19389), .X(n19011) );
  xnor2_1 U19074 ( .A(n11554), .B(n19479), .Y(n19389) );
  nor2_1 U19075 ( .A(outData[4]), .B(outData[6]), .Y(n19479) );
  nand2_1 U19076 ( .A(n19480), .B(n19390), .Y(n19478) );
  nand2_1 U19077 ( .A(n19481), .B(n18593), .Y(n19390) );
  xor2_1 U19078 ( .A(n13368), .B(n19482), .X(n19481) );
  inv_1 U19079 ( .A(n19388), .Y(n19480) );
  nor2_1 U19080 ( .A(n18593), .B(n19483), .Y(n19388) );
  xor2_1 U19081 ( .A(n13351), .B(n19484), .X(n19483) );
  inv_1 U19082 ( .A(n13368), .Y(n13351) );
  xnor2_1 U19083 ( .A(n19485), .B(n19486), .Y(n18593) );
  xor2_1 U19084 ( .A(n18213), .B(n19487), .X(n19485) );
  a21oi_1 U19085 ( .A1(n19488), .A2(n23995), .B1(n19489), .Y(n19487) );
  inv_1 U19086 ( .A(n19490), .Y(n19488) );
  o21ai_0 U19087 ( .A1(n19491), .A2(n19492), .B1(n19493), .Y(n19490) );
  inv_1 U19088 ( .A(n19010), .Y(n19391) );
  nand2_1 U19089 ( .A(n19494), .B(n19418), .Y(n19010) );
  nand2_1 U19090 ( .A(n19495), .B(n18600), .Y(n19418) );
  xor2_1 U19091 ( .A(n18840), .B(n19496), .X(n19495) );
  xor2_1 U19092 ( .A(n17550), .B(n19497), .X(n19494) );
  nand2_1 U19093 ( .A(n19498), .B(n19417), .Y(n19497) );
  o21ai_0 U19094 ( .A1(outData[6]), .A2(n10604), .B1(n19499), .Y(n19417) );
  xor2_1 U19095 ( .A(n18213), .B(n19419), .X(n19498) );
  nand2_1 U19096 ( .A(n19500), .B(n19501), .Y(n19419) );
  inv_1 U19097 ( .A(n18600), .Y(n19501) );
  xnor2_1 U19098 ( .A(n19502), .B(n19503), .Y(n18600) );
  o21ai_0 U19099 ( .A1(n19504), .A2(n19505), .B1(n19506), .Y(n19502) );
  xor2_1 U19100 ( .A(n19496), .B(n19507), .X(n19500) );
  xor2_1 U19101 ( .A(n19508), .B(n12533), .X(n18993) );
  inv_1 U19102 ( .A(n18994), .Y(n18987) );
  o21ai_0 U19103 ( .A1(n19387), .A2(n19509), .B1(n19510), .Y(n18994) );
  mux2i_1 U19104 ( .A0(n19511), .A1(n19512), .S(n12806), .Y(n19510) );
  nor2_1 U19105 ( .A(n19513), .B(n18615), .Y(n19512) );
  mux2i_1 U19106 ( .A0(n19514), .A1(n19515), .S(n16750), .Y(n19509) );
  or2_0 U19107 ( .A(n17240), .B(n19516), .X(n19515) );
  nor2_1 U19108 ( .A(n19513), .B(n17240), .Y(n19514) );
  inv_1 U19109 ( .A(n19386), .Y(n19513) );
  o21ai_0 U19110 ( .A1(n19516), .A2(n17240), .B1(n19511), .Y(n19386) );
  nand2_1 U19111 ( .A(n19516), .B(n17240), .Y(n19511) );
  inv_1 U19112 ( .A(n18615), .Y(n17240) );
  xor2_1 U19113 ( .A(n19517), .B(n19518), .X(n18615) );
  nand2_1 U19114 ( .A(n19519), .B(n19520), .Y(n19517) );
  nand2_1 U19115 ( .A(n19521), .B(n19522), .Y(n19055) );
  o21ai_0 U19116 ( .A1(n19523), .A2(n18582), .B1(n12533), .Y(n19522) );
  mux2i_1 U19117 ( .A0(n19508), .A1(n19524), .S(n13009), .Y(n19521) );
  and2_0 U19118 ( .A(n18582), .B(n19523), .X(n19524) );
  xor2_1 U19119 ( .A(n19523), .B(n18582), .X(n19508) );
  inv_1 U19120 ( .A(n18583), .Y(n18582) );
  xor2_1 U19121 ( .A(n19525), .B(n19526), .X(n18583) );
  xor2_1 U19122 ( .A(n19527), .B(n17391), .X(n19525) );
  inv_1 U19123 ( .A(n16753), .Y(n17391) );
  o221ai_1 U19124 ( .A1(n19528), .A2(n12356), .B1(n19529), .B2(n12411), .C1(
        n19530), .Y(n16753) );
  inv_1 U19125 ( .A(n19531), .Y(n12411) );
  nand2_1 U19126 ( .A(n19532), .B(n19533), .Y(n19527) );
  xnor2_1 U19127 ( .A(n17992), .B(n19534), .Y(n19523) );
  nor2_1 U19128 ( .A(outData[6]), .B(outData[8]), .Y(n19534) );
  xnor2_1 U19129 ( .A(n12789), .B(n19535), .Y(n19053) );
  xor2_1 U19130 ( .A(n18134), .B(n19536), .X(n19535) );
  xor2_1 U19131 ( .A(n17697), .B(n19537), .X(n19377) );
  nor2_1 U19132 ( .A(n18976), .B(n18978), .Y(n19537) );
  xnor2_1 U19133 ( .A(n18576), .B(n19538), .Y(n18976) );
  nor2_1 U19134 ( .A(n19539), .B(n19540), .Y(n19538) );
  o22ai_1 U19135 ( .A1(n19541), .A2(n12789), .B1(n19542), .B2(n18134), .Y(
        n18978) );
  nor2_1 U19136 ( .A(n19536), .B(n19543), .Y(n19542) );
  inv_1 U19137 ( .A(n12789), .Y(n19543) );
  xnor2_1 U19138 ( .A(n19544), .B(n19545), .Y(n12789) );
  xor2_1 U19139 ( .A(n19546), .B(n19547), .X(n19544) );
  xor2_1 U19140 ( .A(n18379), .B(n19548), .X(n19372) );
  nor2_1 U19141 ( .A(n19067), .B(n19068), .Y(n19548) );
  xor2_1 U19142 ( .A(n19549), .B(n19550), .X(n19068) );
  xor2_1 U19143 ( .A(n19551), .B(n18565), .X(n19549) );
  xnor2_1 U19144 ( .A(n17403), .B(n19552), .Y(n19067) );
  a21oi_1 U19145 ( .A1(n18576), .A2(n19553), .B1(n19540), .Y(n19552) );
  and2_0 U19146 ( .A(n19554), .B(n19555), .X(n19540) );
  inv_1 U19147 ( .A(n19539), .Y(n19553) );
  nor2_1 U19148 ( .A(n19555), .B(n19554), .Y(n19539) );
  nand2_1 U19149 ( .A(n12402), .B(n12330), .Y(n19555) );
  xor2_1 U19150 ( .A(n19556), .B(n19557), .X(n18576) );
  nor2_1 U19151 ( .A(n19558), .B(n19559), .Y(n19557) );
  o221ai_1 U19152 ( .A1(n13396), .A2(n13369), .B1(n13383), .B2(n19560), .C1(
        n19561), .Y(n17403) );
  nand2_1 U19153 ( .A(n13397), .B(n24021), .Y(n19561) );
  nor2_1 U19154 ( .A(n13409), .B(n19562), .Y(n13396) );
  xor2_1 U19155 ( .A(n19563), .B(n18559), .X(n19370) );
  xnor2_1 U19156 ( .A(n19564), .B(n19565), .Y(n19563) );
  inv_1 U19157 ( .A(n19077), .Y(n19369) );
  o21ai_0 U19158 ( .A1(n19566), .A2(n19551), .B1(n19567), .Y(n19077) );
  xnor2_1 U19159 ( .A(n11103), .B(n19568), .Y(n19567) );
  nand2_1 U19160 ( .A(n19550), .B(n19569), .Y(n19568) );
  xor2_1 U19161 ( .A(n23995), .B(n19570), .X(n19569) );
  nor2_1 U19162 ( .A(n19571), .B(n18565), .Y(n19570) );
  inv_1 U19163 ( .A(n19566), .Y(n18565) );
  inv_1 U19164 ( .A(n19551), .Y(n19571) );
  nand2_1 U19165 ( .A(n12414), .B(n10611), .Y(n19551) );
  o21ai_0 U19166 ( .A1(n19572), .A2(n19573), .B1(n19574), .Y(n19566) );
  mux2i_1 U19167 ( .A0(n19575), .A1(n19576), .S(n19577), .Y(n19574) );
  nor2_1 U19168 ( .A(n19578), .B(n19503), .Y(n19575) );
  xnor2_1 U19169 ( .A(n19577), .B(n19503), .Y(n19573) );
  or2_0 U19170 ( .A(n19367), .B(n19366), .X(n19084) );
  inv_1 U19171 ( .A(n19579), .Y(n19366) );
  o22ai_1 U19172 ( .A1(n19565), .A2(n18559), .B1(n19564), .B2(n19580), .Y(
        n19579) );
  and2_0 U19173 ( .A(n18559), .B(n19565), .X(n19580) );
  inv_1 U19174 ( .A(n19581), .Y(n18559) );
  o21ai_0 U19175 ( .A1(n19582), .A2(n19583), .B1(n19584), .Y(n19581) );
  mux2i_1 U19176 ( .A0(n19585), .A1(n19586), .S(n19587), .Y(n19584) );
  o21ai_0 U19177 ( .A1(n19588), .A2(n19589), .B1(n19590), .Y(n19585) );
  xor2_1 U19178 ( .A(n24045), .B(n19591), .X(n19590) );
  xor2_1 U19179 ( .A(n19492), .B(n19588), .X(n19583) );
  nor2_1 U19180 ( .A(outData[10]), .B(outData[12]), .Y(n19565) );
  xnor2_1 U19181 ( .A(n18555), .B(n19592), .Y(n19367) );
  a21oi_1 U19182 ( .A1(n19363), .A2(n19593), .B1(n19364), .Y(n19592) );
  nor2_1 U19183 ( .A(n19593), .B(n19363), .Y(n19364) );
  inv_1 U19184 ( .A(n19358), .Y(n18555) );
  xor2_1 U19185 ( .A(n19594), .B(n19595), .X(n19358) );
  nor2_1 U19186 ( .A(n19596), .B(n19597), .Y(n19595) );
  xnor2_1 U19187 ( .A(n19598), .B(n12489), .Y(n19090) );
  xor2_1 U19188 ( .A(n19599), .B(n19600), .X(n19598) );
  inv_1 U19189 ( .A(n18956), .Y(n19351) );
  xor2_1 U19190 ( .A(n19601), .B(n19602), .X(n18956) );
  xor2_1 U19191 ( .A(n19603), .B(n11510), .X(n19602) );
  inv_1 U19192 ( .A(n12956), .Y(n11510) );
  o21ai_0 U19193 ( .A1(n24042), .A2(n14697), .B1(n14666), .Y(n12956) );
  xor2_1 U19194 ( .A(n12529), .B(n19604), .X(n19601) );
  inv_1 U19195 ( .A(n19354), .Y(n18957) );
  o22ai_1 U19196 ( .A1(n19600), .A2(n12489), .B1(n19605), .B2(n19606), .Y(
        n19354) );
  nor2_1 U19197 ( .A(n18132), .B(n19607), .Y(n19606) );
  inv_1 U19198 ( .A(n19607), .Y(n12489) );
  o221ai_1 U19199 ( .A1(n19608), .A2(n19609), .B1(n19610), .B2(n19611), .C1(
        n19612), .Y(n19607) );
  a21oi_1 U19200 ( .A1(n19613), .A2(n19614), .B1(n19615), .Y(n19610) );
  xor2_1 U19201 ( .A(n11684), .B(n19616), .X(n19615) );
  xor2_1 U19202 ( .A(n19617), .B(n19613), .X(n19609) );
  inv_1 U19203 ( .A(n18132), .Y(n19600) );
  xor2_1 U19204 ( .A(n19618), .B(n16868), .X(n19348) );
  nand2_1 U19205 ( .A(n18944), .B(n18943), .Y(n19618) );
  xor2_1 U19206 ( .A(n19619), .B(n19620), .X(n18943) );
  xor2_1 U19207 ( .A(n12543), .B(n19621), .X(n19620) );
  xor2_1 U19208 ( .A(n16845), .B(n16275), .X(n19621) );
  xnor2_1 U19209 ( .A(n18635), .B(n19622), .Y(n19619) );
  inv_1 U19210 ( .A(n19623), .Y(n18944) );
  o22ai_1 U19211 ( .A1(n19624), .A2(n18541), .B1(n19603), .B2(n19625), .Y(
        n19623) );
  nor2_1 U19212 ( .A(n12529), .B(n19604), .Y(n19625) );
  inv_1 U19213 ( .A(n12529), .Y(n18541) );
  xnor2_1 U19214 ( .A(n19626), .B(n19545), .Y(n12529) );
  xor2_1 U19215 ( .A(n19627), .B(n19628), .X(n19626) );
  inv_1 U19216 ( .A(n19604), .Y(n19624) );
  o22ai_1 U19217 ( .A1(n19622), .A2(n18635), .B1(n19629), .B2(n19630), .Y(
        n18937) );
  and2_0 U19218 ( .A(n18635), .B(n19622), .X(n19629) );
  mux2i_1 U19219 ( .A0(n19631), .A1(n19632), .S(n19633), .Y(n18635) );
  xor2_1 U19220 ( .A(n19634), .B(n19635), .X(n19632) );
  xor2_1 U19221 ( .A(n19636), .B(n19635), .X(n19631) );
  xor2_1 U19222 ( .A(n18521), .B(n19637), .X(n19635) );
  xnor2_1 U19223 ( .A(n19638), .B(n16904), .Y(n19622) );
  nand2_1 U19224 ( .A(n12310), .B(n19639), .Y(n19638) );
  xor2_1 U19225 ( .A(n19640), .B(n19641), .X(n18934) );
  xor2_1 U19226 ( .A(n19466), .B(n18642), .X(n19641) );
  o221ai_1 U19227 ( .A1(n19642), .A2(n19643), .B1(n19644), .B2(n19645), .C1(
        n19646), .Y(n18642) );
  a21oi_1 U19228 ( .A1(n19572), .A2(n19647), .B1(n19648), .Y(n19645) );
  xor2_1 U19229 ( .A(n11185), .B(n19649), .X(n19648) );
  xor2_1 U19230 ( .A(n19572), .B(n19650), .X(n19643) );
  xnor2_1 U19231 ( .A(n19334), .B(n19336), .Y(n19640) );
  nor2_1 U19232 ( .A(outData[17]), .B(outData[15]), .Y(n19334) );
  xnor2_1 U19233 ( .A(n12297), .B(n19651), .Y(n19119) );
  a21oi_1 U19234 ( .A1(n19312), .A2(n18525), .B1(n19652), .Y(n19651) );
  xor2_1 U19235 ( .A(n11621), .B(n19653), .X(n19652) );
  nand2_1 U19236 ( .A(n19320), .B(n19654), .Y(n19653) );
  xor2_1 U19237 ( .A(n17715), .B(n19655), .X(n19654) );
  nor2_1 U19238 ( .A(n19312), .B(n18525), .Y(n19655) );
  xor2_1 U19239 ( .A(n10893), .B(n19656), .X(n19320) );
  mux2_1 U19240 ( .A0(n19657), .A1(n19658), .S(n19659), .X(n18525) );
  xor2_1 U19241 ( .A(n19660), .B(n19661), .X(n19658) );
  xor2_1 U19242 ( .A(n19662), .B(n19661), .X(n19657) );
  xor2_1 U19243 ( .A(n17774), .B(n19663), .X(n19661) );
  o22ai_1 U19244 ( .A1(n18508), .A2(n19664), .B1(n19665), .B2(n19297), .Y(
        n19130) );
  xor2_1 U19245 ( .A(n17475), .B(n19666), .X(n19297) );
  inv_1 U19246 ( .A(n18732), .Y(n17475) );
  nand3_1 U19247 ( .A(n19667), .B(n19668), .C(n19669), .Y(n18732) );
  a22oi_1 U19248 ( .A1(n24046), .A2(n19670), .B1(n14650), .B2(n19671), .Y(
        n19669) );
  inv_1 U19249 ( .A(n14702), .Y(n14650) );
  o22ai_1 U19250 ( .A1(n24017), .A2(n14707), .B1(n19671), .B2(n14687), .Y(
        n19670) );
  o21ai_0 U19251 ( .A1(n19146), .A2(n19672), .B1(n14682), .Y(n19667) );
  nor2_1 U19252 ( .A(n19298), .B(n12536), .Y(n19665) );
  inv_1 U19253 ( .A(n18508), .Y(n12536) );
  inv_1 U19254 ( .A(n19664), .Y(n19298) );
  xor2_1 U19255 ( .A(n13010), .B(n19673), .X(n19664) );
  nor2_1 U19256 ( .A(outData[19]), .B(outData[21]), .Y(n19673) );
  xor2_1 U19257 ( .A(n19674), .B(n19675), .X(n18508) );
  nor2_1 U19258 ( .A(n19676), .B(n19677), .Y(n19675) );
  inv_1 U19259 ( .A(n19678), .Y(n19676) );
  xnor2_1 U19260 ( .A(n19679), .B(n19680), .Y(n19131) );
  xnor2_1 U19261 ( .A(n19284), .B(n19681), .Y(n19680) );
  xor2_1 U19262 ( .A(n13410), .B(n17830), .X(n19681) );
  xor2_1 U19263 ( .A(n11223), .B(n19282), .X(n19679) );
  xnor2_1 U19264 ( .A(n19682), .B(n10840), .Y(n19282) );
  nor4_1 U19265 ( .A(n19683), .B(n12298), .C(n19684), .D(n19685), .Y(n10840)
         );
  or2_0 U19266 ( .A(n12301), .B(n12377), .X(n19685) );
  nor2_1 U19267 ( .A(n12409), .B(n24023), .Y(n12377) );
  inv_1 U19268 ( .A(n11844), .Y(n12301) );
  nand3_1 U19269 ( .A(n24035), .B(n12383), .C(n12222), .Y(n11844) );
  nor2_1 U19270 ( .A(n18874), .B(n12403), .Y(n12298) );
  nand2_1 U19271 ( .A(n12426), .B(n17676), .Y(n19682) );
  xor2_1 U19272 ( .A(n19686), .B(n19687), .X(n11223) );
  mux2i_1 U19273 ( .A0(n19688), .A1(n19689), .S(n18077), .Y(n19687) );
  mux2i_1 U19274 ( .A0(n19690), .A1(n19691), .S(n19692), .Y(n19689) );
  a21oi_1 U19275 ( .A1(n19693), .A2(n19636), .B1(n19694), .Y(n19688) );
  a21oi_1 U19276 ( .A1(n19288), .A2(n18505), .B1(n19287), .Y(n18901) );
  nor2_1 U19277 ( .A(n19695), .B(n19696), .Y(n19287) );
  xor2_1 U19278 ( .A(n19650), .B(n19697), .X(n18505) );
  xor2_1 U19279 ( .A(n19698), .B(n19699), .X(n19697) );
  nand2_1 U19280 ( .A(n19696), .B(n19695), .Y(n19288) );
  xnor2_1 U19281 ( .A(n17047), .B(n19700), .Y(n18903) );
  a21oi_1 U19282 ( .A1(n19277), .A2(n19701), .B1(n19273), .Y(n19700) );
  nor3_1 U19283 ( .A(outData[22]), .B(outData[24]), .C(n19277), .Y(n19273) );
  nand2_1 U19284 ( .A(n12426), .B(n17709), .Y(n19701) );
  xnor2_1 U19285 ( .A(n19702), .B(n19703), .Y(n17047) );
  xor2_1 U19286 ( .A(n11574), .B(n19704), .X(n19702) );
  a21oi_1 U19287 ( .A1(n19705), .A2(n13009), .B1(n19706), .Y(n19704) );
  inv_1 U19288 ( .A(n19707), .Y(n19705) );
  o21ai_0 U19289 ( .A1(n19222), .A2(n19343), .B1(n19708), .Y(n19707) );
  xor2_1 U19290 ( .A(n19375), .B(n19709), .X(n19265) );
  nor2_1 U19291 ( .A(n19158), .B(n19165), .Y(n19709) );
  inv_1 U19292 ( .A(n19266), .Y(n19165) );
  a21oi_1 U19293 ( .A1(n19270), .A2(n12944), .B1(n19272), .Y(n19266) );
  nor3_1 U19294 ( .A(outData[23]), .B(outData[25]), .C(n18501), .Y(n19272) );
  o21ai_0 U19295 ( .A1(outData[25]), .A2(outData[23]), .B1(n18501), .Y(n19270)
         );
  xor2_1 U19296 ( .A(n19710), .B(n19711), .X(n18501) );
  nor2_1 U19297 ( .A(n19712), .B(n19713), .Y(n19711) );
  inv_1 U19298 ( .A(n19714), .Y(n19712) );
  xor2_1 U19299 ( .A(n19715), .B(n19716), .X(n19158) );
  xor2_1 U19300 ( .A(n16627), .B(n19717), .X(n19716) );
  xor2_1 U19301 ( .A(n19718), .B(n11734), .X(n19715) );
  inv_1 U19302 ( .A(n12972), .Y(n11734) );
  mux2i_1 U19303 ( .A0(n10624), .A1(n19719), .S(n23972), .Y(n12972) );
  o21ai_0 U19304 ( .A1(n13944), .A2(n10624), .B1(n18668), .Y(n19719) );
  xor2_1 U19305 ( .A(n12968), .B(n19720), .X(n19263) );
  nor2_1 U19306 ( .A(n18879), .B(n18877), .Y(n19720) );
  xnor2_1 U19307 ( .A(n19721), .B(n11284), .Y(n18879) );
  inv_1 U19308 ( .A(n11622), .Y(n11284) );
  mux2i_1 U19309 ( .A0(n19722), .A1(n19723), .S(n11751), .Y(n19721) );
  o22ai_1 U19310 ( .A1(n19724), .A2(n18498), .B1(n19725), .B2(n19726), .Y(
        n19723) );
  and2_0 U19311 ( .A(n18498), .B(n19724), .X(n19726) );
  inv_1 U19312 ( .A(n19717), .Y(n19725) );
  inv_1 U19313 ( .A(n11466), .Y(n18498) );
  nor2_1 U19314 ( .A(n19718), .B(n19717), .Y(n19722) );
  xor2_1 U19315 ( .A(n11466), .B(n19724), .X(n19718) );
  nor2_1 U19316 ( .A(outData[26]), .B(outData[24]), .Y(n19724) );
  xor2_1 U19317 ( .A(n19727), .B(n19728), .X(n11466) );
  xor2_1 U19318 ( .A(n12968), .B(n19729), .X(n19728) );
  o21ai_0 U19319 ( .A1(n19730), .A2(n19731), .B1(n19732), .Y(n19729) );
  inv_1 U19320 ( .A(n19733), .Y(n19732) );
  xnor2_1 U19321 ( .A(n19734), .B(n19735), .Y(n18877) );
  xor2_1 U19322 ( .A(n11205), .B(n19259), .X(n19735) );
  xor2_1 U19323 ( .A(n19257), .B(n19258), .X(n19734) );
  xor2_1 U19324 ( .A(n19736), .B(n19737), .X(n19257) );
  xor2_1 U19325 ( .A(n18801), .B(n19738), .X(n19737) );
  nor2_1 U19326 ( .A(n19171), .B(n19173), .Y(n19242) );
  nand2_1 U19327 ( .A(n19739), .B(n19740), .Y(n19173) );
  o21ai_0 U19328 ( .A1(n19741), .A2(n19742), .B1(n12938), .Y(n19740) );
  xor2_1 U19329 ( .A(n18128), .B(n19251), .X(n19742) );
  mux2i_1 U19330 ( .A0(n19743), .A1(n19253), .S(n18128), .Y(n19739) );
  inv_1 U19331 ( .A(n16763), .Y(n18128) );
  nand3_1 U19332 ( .A(n19744), .B(n19745), .C(n19746), .Y(n16763) );
  a211oi_1 U19333 ( .A1(n19747), .A2(n13821), .B1(n19238), .C1(n13952), .Y(
        n19746) );
  nor2_1 U19334 ( .A(n19253), .B(n12938), .Y(n19743) );
  xor2_1 U19335 ( .A(n19748), .B(n19749), .X(n12938) );
  xor2_1 U19336 ( .A(n18774), .B(n19692), .X(n19749) );
  xor2_1 U19337 ( .A(n19750), .B(n16823), .X(n19748) );
  inv_1 U19338 ( .A(n11336), .Y(n16823) );
  o21ai_0 U19339 ( .A1(n19562), .A2(n13369), .B1(n13402), .Y(n11336) );
  nor2_1 U19340 ( .A(n19252), .B(n19251), .Y(n19253) );
  xor2_1 U19341 ( .A(n19751), .B(n11681), .X(n19171) );
  or2_0 U19342 ( .A(n19231), .B(n19233), .X(n19751) );
  and2_0 U19343 ( .A(n19752), .B(n11411), .X(n19233) );
  nor2_1 U19344 ( .A(n11411), .B(n19752), .Y(n19231) );
  xor2_1 U19345 ( .A(n16535), .B(n19753), .X(n19752) );
  nor2_1 U19346 ( .A(outData[29]), .B(outData[27]), .Y(n19753) );
  o21ai_0 U19347 ( .A1(n19754), .A2(n19226), .B1(n19755), .Y(n11411) );
  mux2i_1 U19348 ( .A0(n19229), .A1(n19756), .S(n19230), .Y(n19755) );
  nor2_1 U19349 ( .A(n18779), .B(n19699), .Y(n19756) );
  inv_1 U19350 ( .A(n19226), .Y(n19699) );
  and2_0 U19351 ( .A(n19226), .B(n18779), .X(n19229) );
  xor2_1 U19352 ( .A(n19230), .B(n18779), .X(n19754) );
  xnor2_1 U19353 ( .A(n19224), .B(n19194), .Y(n18779) );
  xor2_1 U19354 ( .A(outData[29]), .B(outData[31]), .X(n19194) );
  o22ai_1 U19355 ( .A1(n19757), .A2(n10612), .B1(outData[30]), .B2(n19758), 
        .Y(n19224) );
  nor2_1 U19356 ( .A(outData[28]), .B(n19759), .Y(n19758) );
  inv_1 U19357 ( .A(n19759), .Y(n19757) );
  o22ai_1 U19358 ( .A1(n19760), .A2(n18774), .B1(n19761), .B2(n19692), .Y(
        n19230) );
  and2_0 U19359 ( .A(n18774), .B(n19760), .X(n19761) );
  xor2_1 U19360 ( .A(n19762), .B(n11681), .X(n18774) );
  o21ai_0 U19361 ( .A1(n11746), .A2(n10612), .B1(n19195), .Y(n11681) );
  nand2_1 U19362 ( .A(n10612), .B(n11746), .Y(n19195) );
  inv_1 U19363 ( .A(outData[30]), .Y(n11746) );
  xor2_1 U19364 ( .A(n19759), .B(n16880), .X(n19762) );
  o22ai_1 U19365 ( .A1(n12412), .A2(n19763), .B1(outData[29]), .B2(n19764), 
        .Y(n19759) );
  and2_0 U19366 ( .A(n12412), .B(n19763), .X(n19764) );
  inv_1 U19367 ( .A(n19750), .Y(n19760) );
  o22ai_1 U19368 ( .A1(n19765), .A2(n18797), .B1(n19766), .B2(n19738), .Y(
        n19750) );
  nor2_1 U19369 ( .A(n18801), .B(n19736), .Y(n19766) );
  inv_1 U19370 ( .A(n18801), .Y(n18797) );
  xor2_1 U19371 ( .A(n19767), .B(n11048), .X(n18801) );
  xor2_1 U19372 ( .A(n19763), .B(n19251), .X(n19767) );
  xnor2_1 U19373 ( .A(n11498), .B(n12412), .Y(n19251) );
  inv_1 U19374 ( .A(outData[29]), .Y(n11498) );
  o22ai_1 U19375 ( .A1(outData[26]), .A2(n19768), .B1(n19769), .B2(n10612), 
        .Y(n19763) );
  nor2_1 U19376 ( .A(n19770), .B(n17711), .Y(n19769) );
  inv_1 U19377 ( .A(n19770), .Y(n19768) );
  inv_1 U19378 ( .A(n19736), .Y(n19765) );
  xor2_1 U19379 ( .A(n18086), .B(n19771), .X(n19736) );
  a21oi_1 U19380 ( .A1(n19727), .A2(n19772), .B1(n19733), .Y(n19771) );
  nor2_1 U19381 ( .A(n19773), .B(n18811), .Y(n19733) );
  xor2_1 U19382 ( .A(n19730), .B(n17958), .X(n18811) );
  or2_0 U19383 ( .A(n19731), .B(n19730), .X(n19772) );
  xnor2_1 U19384 ( .A(n19770), .B(n19774), .Y(n19730) );
  xor2_1 U19385 ( .A(n11650), .B(n19258), .X(n19774) );
  a21oi_1 U19386 ( .A1(outData[26]), .A2(outData[28]), .B1(n19741), .Y(n19258)
         );
  inv_1 U19387 ( .A(n19252), .Y(n19741) );
  nand2_1 U19388 ( .A(n17711), .B(n10612), .Y(n19252) );
  mux2i_1 U19389 ( .A0(n19775), .A1(n19776), .S(n18563), .Y(n19770) );
  inv_1 U19390 ( .A(n16934), .Y(n18563) );
  o22ai_1 U19391 ( .A1(n11416), .A2(n19777), .B1(outData[27]), .B2(n19778), 
        .Y(n19776) );
  nor2_1 U19392 ( .A(n19779), .B(outData[25]), .Y(n19778) );
  inv_1 U19393 ( .A(n12412), .Y(outData[27]) );
  inv_1 U19394 ( .A(n19779), .Y(n19777) );
  nand2_1 U19395 ( .A(n19779), .B(n19717), .Y(n19775) );
  o21ai_0 U19396 ( .A1(n19713), .A2(n19710), .B1(n19714), .Y(n19727) );
  nand2_1 U19397 ( .A(n19780), .B(n19207), .Y(n19714) );
  o21ai_0 U19398 ( .A1(n19706), .A2(n19708), .B1(n19781), .Y(n19710) );
  o22ai_1 U19399 ( .A1(n19343), .A2(n19222), .B1(n19782), .B2(n19703), .Y(
        n19781) );
  o22ai_1 U19400 ( .A1(n19226), .A2(n19698), .B1(n19783), .B2(n19650), .Y(
        n19703) );
  and2_0 U19401 ( .A(n19698), .B(n19226), .X(n19783) );
  o21ai_0 U19402 ( .A1(n19690), .A2(n19692), .B1(n19784), .Y(n19698) );
  xor2_1 U19403 ( .A(n24045), .B(n19785), .X(n19784) );
  nor2_1 U19404 ( .A(n19694), .B(n19686), .Y(n19785) );
  xor2_1 U19405 ( .A(n12968), .B(n19786), .X(n19686) );
  a21oi_1 U19406 ( .A1(n19674), .A2(n19678), .B1(n19677), .Y(n19786) );
  xor2_1 U19407 ( .A(n12649), .B(n19787), .X(n19677) );
  nor2_1 U19408 ( .A(n19627), .B(n19738), .Y(n19787) );
  xor2_1 U19409 ( .A(n19788), .B(n12297), .X(n19738) );
  nand2_1 U19410 ( .A(n19627), .B(n19789), .Y(n19678) );
  inv_1 U19411 ( .A(n19788), .Y(n19789) );
  xor2_1 U19412 ( .A(n19790), .B(n19791), .X(n19788) );
  xor2_1 U19413 ( .A(n16934), .B(n12881), .X(n19791) );
  inv_1 U19414 ( .A(n18136), .Y(n12881) );
  xor2_1 U19415 ( .A(n19792), .B(n19284), .X(n19790) );
  inv_1 U19416 ( .A(n19793), .Y(n19284) );
  a21oi_1 U19417 ( .A1(outData[23]), .A2(outData[21]), .B1(n19696), .Y(n19793)
         );
  nor2_1 U19418 ( .A(outData[23]), .B(outData[21]), .Y(n19696) );
  nand2_1 U19419 ( .A(n19794), .B(n19306), .Y(n19674) );
  xnor2_1 U19420 ( .A(n16275), .B(n19795), .Y(n19306) );
  nor2_1 U19421 ( .A(n19796), .B(n19731), .Y(n19795) );
  xor2_1 U19422 ( .A(n19773), .B(n17765), .X(n19731) );
  xor2_1 U19423 ( .A(n17573), .B(n19797), .X(n19794) );
  nand2_1 U19424 ( .A(n19304), .B(n19305), .Y(n19797) );
  xnor2_1 U19425 ( .A(n11292), .B(n19798), .Y(n19305) );
  nor2_1 U19426 ( .A(n19617), .B(n19773), .Y(n19798) );
  xnor2_1 U19427 ( .A(n19799), .B(n19666), .Y(n19773) );
  xor2_1 U19428 ( .A(outData[20]), .B(n12426), .X(n19666) );
  xor2_1 U19429 ( .A(n19800), .B(n19453), .X(n19799) );
  inv_1 U19430 ( .A(n16666), .Y(n19453) );
  xnor2_1 U19431 ( .A(n19801), .B(n13368), .Y(n19304) );
  o22ai_1 U19432 ( .A1(n19660), .A2(n19663), .B1(n19802), .B2(n19659), .Y(
        n19801) );
  inv_1 U19433 ( .A(n19803), .Y(n19659) );
  and2_0 U19434 ( .A(n19663), .B(n19780), .X(n19802) );
  o22ai_1 U19435 ( .A1(n19345), .A2(n19344), .B1(n19804), .B2(n19343), .Y(
        n19663) );
  and2_0 U19436 ( .A(n19344), .B(n19588), .X(n19804) );
  o221ai_1 U19437 ( .A1(n19649), .A2(n19642), .B1(n19650), .B2(n19578), .C1(
        n19646), .Y(n19344) );
  nand3_1 U19438 ( .A(n19644), .B(n11185), .C(n19649), .Y(n19646) );
  inv_1 U19439 ( .A(n17715), .Y(n11185) );
  inv_1 U19440 ( .A(n19647), .Y(n19650) );
  nand2_1 U19441 ( .A(n19644), .B(n17715), .Y(n19642) );
  a221oi_1 U19442 ( .A1(n14671), .A2(n14596), .B1(n14707), .B2(n19672), .C1(
        n19805), .Y(n17715) );
  inv_1 U19443 ( .A(n14663), .Y(n19672) );
  inv_1 U19444 ( .A(n14673), .Y(n14671) );
  inv_1 U19445 ( .A(n19806), .Y(n19644) );
  o22ai_1 U19446 ( .A1(n19634), .A2(n19637), .B1(n19807), .B2(n19633), .Y(
        n19806) );
  and2_0 U19447 ( .A(n19637), .B(n19690), .X(n19807) );
  o22ai_1 U19448 ( .A1(n19628), .A2(n19808), .B1(n19809), .B2(n19545), .Y(
        n19637) );
  nor2_1 U19449 ( .A(n19627), .B(n19810), .Y(n19809) );
  inv_1 U19450 ( .A(n19808), .Y(n19627) );
  xnor2_1 U19451 ( .A(n19630), .B(n19811), .Y(n19808) );
  inv_1 U19452 ( .A(n12543), .Y(n19630) );
  xnor2_1 U19453 ( .A(n17633), .B(n12346), .Y(n12543) );
  inv_1 U19454 ( .A(n19810), .Y(n19628) );
  o221ai_1 U19455 ( .A1(n19616), .A2(n19608), .B1(n19617), .B2(n19812), .C1(
        n19612), .Y(n19810) );
  nand3_1 U19456 ( .A(n19616), .B(n19611), .C(n11684), .Y(n19612) );
  inv_1 U19457 ( .A(n12512), .Y(n11684) );
  nand2_1 U19458 ( .A(n19611), .B(n12512), .Y(n19608) );
  nand2_1 U19459 ( .A(n19813), .B(n19814), .Y(n12512) );
  o211ai_1 U19460 ( .A1(n24007), .A2(n16177), .B1(n16187), .C1(n16190), .Y(
        n19813) );
  o21ai_0 U19461 ( .A1(n19815), .A2(n19596), .B1(n19816), .Y(n19611) );
  inv_1 U19462 ( .A(n19597), .Y(n19816) );
  xor2_1 U19463 ( .A(n19817), .B(n19818), .X(n19597) );
  nor2_1 U19464 ( .A(n19819), .B(n19803), .Y(n19818) );
  xor2_1 U19465 ( .A(n13014), .B(n19820), .X(n19596) );
  and2_0 U19466 ( .A(n19803), .B(n19819), .X(n19820) );
  xnor2_1 U19467 ( .A(n19821), .B(n19605), .Y(n19803) );
  inv_1 U19468 ( .A(n19594), .Y(n19815) );
  o221ai_1 U19469 ( .A1(n19591), .A2(n19582), .B1(n19588), .B2(n19589), .C1(
        n19822), .Y(n19594) );
  nand2_1 U19470 ( .A(n19586), .B(n19587), .Y(n19822) );
  and2_0 U19471 ( .A(n19591), .B(n14685), .X(n19586) );
  inv_1 U19472 ( .A(n19492), .Y(n19589) );
  inv_1 U19473 ( .A(n19346), .Y(n19588) );
  nand2_1 U19474 ( .A(n24045), .B(n19587), .Y(n19582) );
  o21ai_0 U19475 ( .A1(n19572), .A2(n19503), .B1(n19823), .Y(n19587) );
  xor2_1 U19476 ( .A(n18405), .B(n19824), .X(n19823) );
  or2_0 U19477 ( .A(n19577), .B(n19576), .X(n19824) );
  and2_0 U19478 ( .A(n19572), .B(n19503), .X(n19576) );
  xor2_1 U19479 ( .A(n19825), .B(n18204), .X(n19577) );
  inv_1 U19480 ( .A(n13010), .Y(n18204) );
  nand2_1 U19481 ( .A(n19826), .B(n19827), .Y(n19825) );
  inv_1 U19482 ( .A(n19559), .Y(n19827) );
  xor2_1 U19483 ( .A(n18947), .B(n19828), .X(n19559) );
  nor2_1 U19484 ( .A(n19633), .B(n19829), .Y(n19828) );
  xnor2_1 U19485 ( .A(n18521), .B(n19830), .Y(n19826) );
  nor2_1 U19486 ( .A(n19558), .B(n19556), .Y(n19830) );
  o22ai_1 U19487 ( .A1(n19545), .A2(n19547), .B1(n19831), .B2(n19546), .Y(
        n19556) );
  inv_1 U19488 ( .A(n19477), .Y(n19546) );
  and2_0 U19489 ( .A(n19547), .B(n19545), .X(n19831) );
  xnor2_1 U19490 ( .A(n17616), .B(n19832), .Y(n19547) );
  a21oi_1 U19491 ( .A1(n19526), .A2(n19532), .B1(n19833), .Y(n19832) );
  inv_1 U19492 ( .A(n19533), .Y(n19833) );
  nand2_1 U19493 ( .A(n19457), .B(n19812), .Y(n19533) );
  xor2_1 U19494 ( .A(n16995), .B(n19834), .X(n19532) );
  nor2_1 U19495 ( .A(n19457), .B(n19812), .Y(n19834) );
  inv_1 U19496 ( .A(n19613), .Y(n19812) );
  xor2_1 U19497 ( .A(n19835), .B(n18125), .X(n19526) );
  nand2_1 U19498 ( .A(n19836), .B(n19520), .Y(n19835) );
  nand2_1 U19499 ( .A(n19819), .B(n19461), .Y(n19520) );
  xnor2_1 U19500 ( .A(n19837), .B(n19838), .Y(n19836) );
  nand2_1 U19501 ( .A(n19518), .B(n19519), .Y(n19838) );
  or2_0 U19502 ( .A(n19461), .B(n19819), .X(n19519) );
  xor2_1 U19503 ( .A(n12533), .B(n19839), .X(n19819) );
  xor2_1 U19504 ( .A(n19840), .B(n12968), .X(n19518) );
  o22ai_1 U19505 ( .A1(n19492), .A2(n19491), .B1(n19841), .B2(n19486), .Y(
        n19840) );
  xor2_1 U19506 ( .A(n16868), .B(n19842), .X(n19486) );
  and2_0 U19507 ( .A(n19843), .B(n19506), .X(n19842) );
  nand2_1 U19508 ( .A(n19504), .B(n19505), .Y(n19506) );
  o21ai_0 U19509 ( .A1(n19505), .A2(n19504), .B1(n19503), .Y(n19843) );
  a21oi_1 U19510 ( .A1(outData[1]), .A2(outData[0]), .B1(n18138), .Y(n19504)
         );
  o21ai_0 U19511 ( .A1(n12464), .A2(n19468), .B1(n19844), .Y(n19505) );
  xor2_1 U19512 ( .A(n18021), .B(n19845), .X(n19844) );
  a21oi_1 U19513 ( .A1(n19468), .A2(n12464), .B1(n19467), .Y(n19845) );
  nand2_1 U19514 ( .A(n19458), .B(n19477), .Y(n19467) );
  xnor2_1 U19515 ( .A(n19846), .B(n19847), .Y(n19477) );
  nor2_1 U19516 ( .A(n19456), .B(n19457), .Y(n19458) );
  mux2_1 U19517 ( .A0(n19848), .A1(n19849), .S(outData[2]), .X(n19457) );
  inv_1 U19518 ( .A(n12308), .Y(outData[2]) );
  xor2_1 U19519 ( .A(n10604), .B(n19850), .X(n19849) );
  xor2_1 U19520 ( .A(n19851), .B(n19850), .X(n19848) );
  or2_0 U19521 ( .A(n19452), .B(n19461), .X(n19456) );
  xnor2_1 U19522 ( .A(n19440), .B(n19852), .Y(n19461) );
  xor2_1 U19523 ( .A(n10919), .B(n19853), .X(n19852) );
  inv_1 U19524 ( .A(n19443), .Y(n19440) );
  a21oi_1 U19525 ( .A1(outData[1]), .A2(outData[3]), .B1(n19439), .Y(n19443)
         );
  nor2_1 U19526 ( .A(outData[1]), .B(outData[3]), .Y(n19439) );
  inv_1 U19527 ( .A(n12506), .Y(outData[1]) );
  xor2_1 U19528 ( .A(n17578), .B(n17830), .X(n19452) );
  o221ai_1 U19529 ( .A1(n13929), .A2(n13950), .B1(n23990), .B2(n19234), .C1(
        n19854), .Y(n17830) );
  a221oi_1 U19530 ( .A1(n13924), .A2(n13928), .B1(n13885), .B2(n19855), .C1(
        n19856), .Y(n19854) );
  nor2_1 U19531 ( .A(n13928), .B(n23991), .Y(n13885) );
  nand2_1 U19532 ( .A(n18138), .B(n12308), .Y(n17578) );
  inv_1 U19533 ( .A(n19829), .Y(n19468) );
  a21oi_1 U19534 ( .A1(n23995), .A2(n19493), .B1(n19489), .Y(n19841) );
  nor2_1 U19535 ( .A(n19493), .B(n23995), .Y(n19489) );
  nand2_1 U19536 ( .A(n19492), .B(n19491), .Y(n19493) );
  xor2_1 U19537 ( .A(n19449), .B(n19040), .X(n19491) );
  nand3_1 U19538 ( .A(n19857), .B(n19858), .C(n19859), .Y(n17616) );
  nor3_1 U19539 ( .A(n19860), .B(n19861), .C(n12294), .Y(n19859) );
  inv_1 U19540 ( .A(n19862), .Y(n12294) );
  and3_1 U19541 ( .A(n19318), .B(n10610), .C(n12387), .X(n19860) );
  mux2i_1 U19542 ( .A0(n19863), .A1(n19864), .S(n24027), .Y(n19857) );
  or2_0 U19543 ( .A(n12283), .B(n19865), .X(n19863) );
  nor3_1 U19544 ( .A(n12387), .B(n24030), .C(n12374), .Y(n12283) );
  xor2_1 U19545 ( .A(n19554), .B(n19866), .X(n19545) );
  xor2_1 U19546 ( .A(n10611), .B(outData[9]), .X(n19554) );
  and2_0 U19547 ( .A(n19633), .B(n19829), .X(n19558) );
  o21ai_0 U19548 ( .A1(outData[6]), .A2(n19867), .B1(n19868), .Y(n19829) );
  mux2i_1 U19549 ( .A0(n19869), .A1(n19870), .S(n19871), .Y(n19868) );
  inv_1 U19550 ( .A(n19499), .Y(n19870) );
  nor2_1 U19551 ( .A(n10619), .B(n10604), .Y(n19869) );
  xor2_1 U19552 ( .A(n19871), .B(n19851), .X(n19867) );
  xor2_1 U19553 ( .A(n19550), .B(n19872), .X(n19633) );
  xor2_1 U19554 ( .A(outData[12]), .B(outData[10]), .X(n19550) );
  o221ai_1 U19555 ( .A1(n12357), .A2(n12356), .B1(n19528), .B2(n19529), .C1(
        n19873), .Y(n18521) );
  mux2i_1 U19556 ( .A0(n19874), .A1(n19875), .S(n12384), .Y(n19873) );
  nand2_1 U19557 ( .A(n12423), .B(n12425), .Y(n19874) );
  xor2_1 U19558 ( .A(n19876), .B(n19482), .X(n19503) );
  xor2_1 U19559 ( .A(n17133), .B(n19877), .X(n19876) );
  nor2_1 U19560 ( .A(n19346), .B(n19492), .Y(n19591) );
  xor2_1 U19561 ( .A(n19878), .B(n19879), .X(n19492) );
  xor2_1 U19562 ( .A(n17697), .B(n19387), .X(n19879) );
  xor2_1 U19563 ( .A(n10619), .B(outData[8]), .X(n19387) );
  xor2_1 U19564 ( .A(n19345), .B(n18651), .X(n19346) );
  inv_1 U19565 ( .A(n12649), .Y(n18651) );
  o221ai_1 U19566 ( .A1(n12423), .A2(n12356), .B1(n19875), .B2(n19529), .C1(
        n12415), .Y(n12649) );
  nand2_1 U19567 ( .A(n12390), .B(n12406), .Y(n12415) );
  nor2_1 U19568 ( .A(n19614), .B(n19613), .Y(n19616) );
  xor2_1 U19569 ( .A(n19880), .B(n19881), .X(n19613) );
  xor2_1 U19570 ( .A(n11159), .B(n19541), .X(n19880) );
  inv_1 U19571 ( .A(n19536), .Y(n19541) );
  o21ai_0 U19572 ( .A1(n12330), .A2(outData[10]), .B1(n19882), .Y(n19536) );
  inv_1 U19573 ( .A(n19617), .Y(n19614) );
  xor2_1 U19574 ( .A(n19796), .B(n19507), .X(n19617) );
  xor2_1 U19575 ( .A(n19883), .B(n19604), .X(n19796) );
  nor2_1 U19576 ( .A(n19647), .B(n19572), .Y(n19649) );
  inv_1 U19577 ( .A(n19578), .Y(n19572) );
  xor2_1 U19578 ( .A(n19564), .B(n19884), .X(n19578) );
  a21oi_1 U19579 ( .A1(outData[13]), .A2(outData[11]), .B1(n19360), .Y(n19564)
         );
  inv_1 U19580 ( .A(n19593), .Y(n19360) );
  nand2_1 U19581 ( .A(n12413), .B(n10611), .Y(n19593) );
  xnor2_1 U19582 ( .A(n19885), .B(n19324), .Y(n19647) );
  xor2_1 U19583 ( .A(n19886), .B(n19363), .X(n19345) );
  o21ai_0 U19584 ( .A1(n19639), .A2(n10617), .B1(n18132), .Y(n19363) );
  nand2_1 U19585 ( .A(n10617), .B(n19639), .Y(n18132) );
  inv_1 U19586 ( .A(n23903), .Y(n12968) );
  nor2_1 U19587 ( .A(n19691), .B(n19693), .Y(n19694) );
  inv_1 U19588 ( .A(n19692), .Y(n19693) );
  inv_1 U19589 ( .A(n19634), .Y(n19691) );
  xnor2_1 U19590 ( .A(n13410), .B(n19636), .Y(n19634) );
  inv_1 U19591 ( .A(n19690), .Y(n19636) );
  xor2_1 U19592 ( .A(n19887), .B(n19695), .X(n19692) );
  xor2_1 U19593 ( .A(n12426), .B(n17709), .X(n19695) );
  xor2_1 U19594 ( .A(n19336), .B(n19888), .X(n19690) );
  xor2_1 U19595 ( .A(outData[16]), .B(n11225), .X(n19336) );
  xnor2_1 U19596 ( .A(n19889), .B(n19277), .Y(n19226) );
  xnor2_1 U19597 ( .A(outData[23]), .B(outData[25]), .Y(n19277) );
  nor2_1 U19598 ( .A(n13009), .B(n19706), .Y(n19782) );
  nor2_1 U19599 ( .A(n19708), .B(n13009), .Y(n19706) );
  inv_1 U19600 ( .A(n18968), .Y(n13009) );
  o211ai_1 U19601 ( .A1(n19890), .A2(n13960), .B1(n16148), .C1(n19891), .Y(
        n18968) );
  nand2_1 U19602 ( .A(n13868), .B(n13916), .Y(n16148) );
  nand2_1 U19603 ( .A(n19343), .B(n19222), .Y(n19708) );
  inv_1 U19604 ( .A(n19208), .Y(n19222) );
  xor2_1 U19605 ( .A(n19892), .B(n12944), .X(n19208) );
  xnor2_1 U19606 ( .A(n17711), .B(outData[24]), .Y(n12944) );
  xnor2_1 U19607 ( .A(n19656), .B(n19893), .Y(n19343) );
  a21oi_1 U19608 ( .A1(n12297), .A2(n19894), .B1(n19895), .Y(n19893) );
  xor2_1 U19609 ( .A(n17676), .B(n11225), .X(n19656) );
  inv_1 U19610 ( .A(outData[18]), .Y(n11225) );
  xor2_1 U19611 ( .A(n11650), .B(n19896), .X(n19713) );
  nor2_1 U19612 ( .A(n19780), .B(n19207), .Y(n19896) );
  xnor2_1 U19613 ( .A(n19717), .B(n19779), .Y(n19207) );
  a21oi_1 U19614 ( .A1(n17709), .A2(n19897), .B1(n19898), .Y(n19779) );
  a21oi_1 U19615 ( .A1(n19892), .A2(outData[24]), .B1(n17711), .Y(n19898) );
  inv_1 U19616 ( .A(outData[26]), .Y(n17711) );
  inv_1 U19617 ( .A(n19892), .Y(n19897) );
  o22ai_1 U19618 ( .A1(n12391), .A2(n19899), .B1(outData[25]), .B2(n19900), 
        .Y(n19892) );
  nor2_1 U19619 ( .A(outData[23]), .B(n19889), .Y(n19900) );
  inv_1 U19620 ( .A(n19889), .Y(n19899) );
  o22ai_1 U19621 ( .A1(n12426), .A2(n19887), .B1(outData[24]), .B2(n19901), 
        .Y(n19889) );
  nor2_1 U19622 ( .A(outData[22]), .B(n19902), .Y(n19901) );
  inv_1 U19623 ( .A(n19887), .Y(n19902) );
  xor2_1 U19624 ( .A(n19903), .B(n18052), .X(n19887) );
  o22ai_1 U19625 ( .A1(outData[23]), .A2(n19792), .B1(n19904), .B2(n11468), 
        .Y(n19903) );
  nor2_1 U19626 ( .A(n12391), .B(n19905), .Y(n19904) );
  inv_1 U19627 ( .A(n19905), .Y(n19792) );
  o22ai_1 U19628 ( .A1(outData[22]), .A2(n19800), .B1(n19906), .B2(n17676), 
        .Y(n19905) );
  and2_0 U19629 ( .A(n19800), .B(outData[22]), .X(n19906) );
  o22ai_1 U19630 ( .A1(outData[19]), .A2(n19907), .B1(n19908), .B2(n11468), 
        .Y(n19800) );
  inv_1 U19631 ( .A(outData[21]), .Y(n11468) );
  nor2_1 U19632 ( .A(n17051), .B(n19909), .Y(n19908) );
  inv_1 U19633 ( .A(n19907), .Y(n19909) );
  inv_1 U19634 ( .A(n12426), .Y(outData[22]) );
  inv_1 U19635 ( .A(n12391), .Y(outData[23]) );
  inv_1 U19636 ( .A(outData[24]), .Y(n17709) );
  o21ai_0 U19637 ( .A1(n12412), .A2(n11416), .B1(n19259), .Y(n19717) );
  nand2_1 U19638 ( .A(n12412), .B(n11416), .Y(n19259) );
  inv_1 U19639 ( .A(outData[25]), .Y(n11416) );
  inv_1 U19640 ( .A(n19662), .Y(n19780) );
  xor2_1 U19641 ( .A(n19660), .B(n16880), .X(n19662) );
  inv_1 U19642 ( .A(n18184), .Y(n16880) );
  xnor2_1 U19643 ( .A(n19907), .B(n12978), .Y(n19660) );
  xor2_1 U19644 ( .A(outData[19]), .B(outData[21]), .X(n12978) );
  xnor2_1 U19645 ( .A(n19910), .B(n12959), .Y(n19907) );
  o22ai_1 U19646 ( .A1(n24006), .A2(n19911), .B1(n16116), .B2(n16187), .Y(
        n12959) );
  o22ai_1 U19647 ( .A1(outData[18]), .A2(n19912), .B1(n19913), .B2(n17676), 
        .Y(n19910) );
  inv_1 U19648 ( .A(outData[20]), .Y(n17676) );
  and2_0 U19649 ( .A(outData[18]), .B(n19912), .X(n19913) );
  nor2_1 U19650 ( .A(n19895), .B(n19914), .Y(n19912) );
  inv_1 U19651 ( .A(n19894), .Y(n19914) );
  o211ai_1 U19652 ( .A1(n12346), .A2(n19885), .B1(n19915), .C1(n12297), .Y(
        n19894) );
  o21ai_0 U19653 ( .A1(outData[17]), .A2(n19916), .B1(n17051), .Y(n19915) );
  inv_1 U19654 ( .A(outData[19]), .Y(n17051) );
  inv_1 U19655 ( .A(n19885), .Y(n19916) );
  nor3_1 U19656 ( .A(n19324), .B(n12297), .C(n19885), .Y(n19895) );
  xor2_1 U19657 ( .A(n19917), .B(n19241), .X(n19885) );
  o22ai_1 U19658 ( .A1(n12310), .A2(n19888), .B1(outData[18]), .B2(n19918), 
        .Y(n19917) );
  and2_0 U19659 ( .A(n12310), .B(n19888), .X(n19918) );
  o22ai_1 U19660 ( .A1(n12346), .A2(n19811), .B1(outData[15]), .B2(n19919), 
        .Y(n19888) );
  nor2_1 U19661 ( .A(outData[17]), .B(n19920), .Y(n19919) );
  inv_1 U19662 ( .A(n19920), .Y(n19811) );
  mux2i_1 U19663 ( .A0(n19921), .A1(n19922), .S(n17598), .Y(n19920) );
  nand2_1 U19664 ( .A(n19923), .B(n19604), .Y(n19922) );
  xnor2_1 U19665 ( .A(n19639), .B(n12310), .Y(n19604) );
  o22ai_1 U19666 ( .A1(outData[16]), .A2(n19883), .B1(n19924), .B2(n19639), 
        .Y(n19921) );
  inv_1 U19667 ( .A(outData[14]), .Y(n19639) );
  nor2_1 U19668 ( .A(n12310), .B(n19923), .Y(n19924) );
  inv_1 U19669 ( .A(n19883), .Y(n19923) );
  mux2i_1 U19670 ( .A0(n19925), .A1(n19926), .S(n17758), .Y(n19883) );
  inv_1 U19671 ( .A(n13014), .Y(n17758) );
  o221ai_1 U19672 ( .A1(n23998), .A2(n13948), .B1(n13868), .B2(n13960), .C1(
        n19396), .Y(n13014) );
  o22ai_1 U19673 ( .A1(outData[15]), .A2(n19927), .B1(n12413), .B2(n19928), 
        .Y(n19926) );
  nor2_1 U19674 ( .A(n17633), .B(n19821), .Y(n19928) );
  inv_1 U19675 ( .A(outData[15]), .Y(n17633) );
  inv_1 U19676 ( .A(n19821), .Y(n19927) );
  nand2_1 U19677 ( .A(n19821), .B(n19599), .Y(n19925) );
  inv_1 U19678 ( .A(n19605), .Y(n19599) );
  a21oi_1 U19679 ( .A1(outData[13]), .A2(outData[15]), .B1(n19603), .Y(n19605)
         );
  nor2_1 U19680 ( .A(outData[13]), .B(outData[15]), .Y(n19603) );
  inv_1 U19681 ( .A(n12413), .Y(outData[13]) );
  o22ai_1 U19682 ( .A1(n10617), .A2(n19929), .B1(outData[14]), .B2(n19930), 
        .Y(n19821) );
  nor2_1 U19683 ( .A(outData[12]), .B(n19886), .Y(n19930) );
  inv_1 U19684 ( .A(n19886), .Y(n19929) );
  xnor2_1 U19685 ( .A(n19931), .B(n12686), .Y(n19886) );
  o22ai_1 U19686 ( .A1(n12413), .A2(n19884), .B1(outData[11]), .B2(n19932), 
        .Y(n19931) );
  and2_0 U19687 ( .A(n12413), .B(n19884), .X(n19932) );
  a21oi_1 U19688 ( .A1(n12402), .A2(n19872), .B1(n19933), .Y(n19884) );
  inv_1 U19689 ( .A(n19934), .Y(n19933) );
  o21ai_0 U19690 ( .A1(n12402), .A2(n19872), .B1(outData[12]), .Y(n19934) );
  o22ai_1 U19691 ( .A1(outData[9]), .A2(n19935), .B1(n19936), .B2(n10611), .Y(
        n19872) );
  nor2_1 U19692 ( .A(n12414), .B(n19866), .Y(n19936) );
  inv_1 U19693 ( .A(n19866), .Y(n19935) );
  o21ai_0 U19694 ( .A1(n19937), .A2(n19881), .B1(n19882), .Y(n19866) );
  nand2_1 U19695 ( .A(n12330), .B(outData[10]), .Y(n19882) );
  mux2_1 U19696 ( .A0(n19938), .A1(n19939), .S(n17591), .X(n19881) );
  nand2_1 U19697 ( .A(n19940), .B(n12533), .Y(n19939) );
  o21ai_0 U19698 ( .A1(n12414), .A2(n17970), .B1(n18134), .Y(n12533) );
  nand2_1 U19699 ( .A(n12414), .B(n17970), .Y(n18134) );
  o22ai_1 U19700 ( .A1(outData[9]), .A2(n19839), .B1(n19941), .B2(n17970), .Y(
        n19938) );
  nor2_1 U19701 ( .A(n12414), .B(n19940), .Y(n19941) );
  inv_1 U19702 ( .A(n19940), .Y(n19839) );
  o22ai_1 U19703 ( .A1(outData[8]), .A2(n19878), .B1(n19942), .B2(n10619), .Y(
        n19940) );
  and2_0 U19704 ( .A(outData[8]), .B(n19878), .X(n19942) );
  mux2i_1 U19705 ( .A0(n19943), .A1(n19944), .S(n18068), .Y(n19878) );
  o22ai_1 U19706 ( .A1(outData[7]), .A2(n19945), .B1(n12440), .B2(n19946), .Y(
        n19944) );
  nor2_1 U19707 ( .A(n19877), .B(n17970), .Y(n19946) );
  inv_1 U19708 ( .A(outData[7]), .Y(n17970) );
  nand2_1 U19709 ( .A(n19877), .B(n19484), .Y(n19943) );
  inv_1 U19710 ( .A(n19482), .Y(n19484) );
  a21oi_1 U19711 ( .A1(outData[5]), .A2(outData[7]), .B1(n19516), .Y(n19482)
         );
  nor2_1 U19712 ( .A(outData[5]), .B(outData[7]), .Y(n19516) );
  inv_1 U19713 ( .A(n19945), .Y(n19877) );
  nand2_1 U19714 ( .A(n19499), .B(n19947), .Y(n19945) );
  o21ai_0 U19715 ( .A1(outData[6]), .A2(n19948), .B1(n19871), .Y(n19947) );
  mux2i_1 U19716 ( .A0(n19949), .A1(n19950), .S(n16801), .Y(n19871) );
  nand4_1 U19717 ( .A(n19951), .B(n19952), .C(n19953), .D(n19954), .Y(n16801)
         );
  a21oi_1 U19718 ( .A1(n19955), .A2(n23978), .B1(n19956), .Y(n19954) );
  mux2i_1 U19719 ( .A0(n16139), .A1(n16121), .S(n16134), .Y(n19956) );
  nand3_1 U19720 ( .A(n23974), .B(n23975), .C(n16107), .Y(n19953) );
  nand2_1 U19721 ( .A(n19957), .B(n19462), .Y(n19950) );
  inv_1 U19722 ( .A(n19847), .Y(n19462) );
  a21oi_1 U19723 ( .A1(outData[5]), .A2(outData[3]), .B1(n19496), .Y(n19847)
         );
  nor2_1 U19724 ( .A(outData[3]), .B(outData[5]), .Y(n19496) );
  o22ai_1 U19725 ( .A1(n12354), .A2(n19846), .B1(outData[5]), .B2(n19958), .Y(
        n19949) );
  nor2_1 U19726 ( .A(outData[3]), .B(n19957), .Y(n19958) );
  inv_1 U19727 ( .A(n19846), .Y(n19957) );
  inv_1 U19728 ( .A(n12440), .Y(outData[5]) );
  xor2_1 U19729 ( .A(n19959), .B(n18458), .X(n19846) );
  inv_1 U19730 ( .A(n19960), .Y(n18458) );
  o22ai_1 U19731 ( .A1(n19850), .A2(n19851), .B1(n12308), .B2(n19961), .Y(
        n19959) );
  nor2_1 U19732 ( .A(n10604), .B(n19962), .Y(n19961) );
  inv_1 U19733 ( .A(n19948), .Y(n19851) );
  inv_1 U19734 ( .A(n19962), .Y(n19850) );
  o22ai_1 U19735 ( .A1(outData[3]), .A2(n19853), .B1(n12506), .B2(n19963), .Y(
        n19962) );
  and2_0 U19736 ( .A(n19853), .B(outData[3]), .X(n19963) );
  o21ai_0 U19737 ( .A1(n18138), .A2(n19964), .B1(n19965), .Y(n19853) );
  mux2i_1 U19738 ( .A0(n11554), .A1(n19966), .S(n12308), .Y(n19965) );
  nor2_1 U19739 ( .A(n11554), .B(outData[0]), .Y(n19966) );
  inv_1 U19740 ( .A(n19168), .Y(n11554) );
  o221ai_1 U19741 ( .A1(n23998), .A2(n19967), .B1(n19968), .B2(n13947), .C1(
        n19891), .Y(n19168) );
  nand2_1 U19742 ( .A(n13867), .B(n23998), .Y(n19891) );
  inv_1 U19743 ( .A(n19040), .Y(n18138) );
  nand2_1 U19744 ( .A(n12464), .B(n12506), .Y(n19040) );
  inv_1 U19745 ( .A(n12354), .Y(outData[3]) );
  xnor2_1 U19746 ( .A(n10604), .B(n10942), .Y(n19948) );
  inv_1 U19747 ( .A(n19969), .Y(n10942) );
  o21ai_0 U19748 ( .A1(n13868), .A2(n19970), .B1(n19971), .Y(n19969) );
  mux2i_1 U19749 ( .A0(n13916), .A1(n24001), .S(n13915), .Y(n19971) );
  nand2_1 U19750 ( .A(outData[6]), .B(n10604), .Y(n19499) );
  inv_1 U19751 ( .A(n12330), .Y(outData[8]) );
  nor2_1 U19752 ( .A(n12330), .B(outData[10]), .Y(n19937) );
  inv_1 U19753 ( .A(n12402), .Y(outData[10]) );
  inv_1 U19754 ( .A(n12414), .Y(outData[9]) );
  inv_1 U19755 ( .A(n12310), .Y(outData[16]) );
  a21oi_1 U19756 ( .A1(outData[17]), .A2(outData[19]), .B1(n19312), .Y(n19324)
         );
  nor2_1 U19757 ( .A(outData[17]), .B(outData[19]), .Y(n19312) );
  inv_1 U19758 ( .A(n12346), .Y(outData[17]) );
  xor2_1 U19759 ( .A(n19972), .B(n19973), .X(n11639) );
  xor2_1 U19760 ( .A(n17598), .B(n19974), .X(n19973) );
  xor2_1 U19761 ( .A(n17000), .B(n24045), .X(n19974) );
  xor2_1 U19762 ( .A(n19975), .B(n16314), .X(n19972) );
  xor2_1 U19763 ( .A(n19976), .B(n18766), .X(n18760) );
  o22ai_1 U19764 ( .A1(n18821), .A2(n11755), .B1(n19977), .B2(n10737), .Y(
        n18766) );
  inv_1 U19765 ( .A(n12476), .Y(n10737) );
  nor2_1 U19766 ( .A(n16730), .B(n19978), .Y(n19977) );
  inv_1 U19767 ( .A(n11755), .Y(n16730) );
  xor2_1 U19768 ( .A(n19979), .B(n19980), .X(n11755) );
  and2_0 U19769 ( .A(n19981), .B(n19982), .X(n19980) );
  xor2_1 U19770 ( .A(n19983), .B(n23903), .X(n19979) );
  nand2_1 U19771 ( .A(n19984), .B(n19985), .Y(n19983) );
  inv_1 U19772 ( .A(n19978), .Y(n18821) );
  o21ai_0 U19773 ( .A1(n18828), .A2(n18826), .B1(n19986), .Y(n19978) );
  inv_1 U19774 ( .A(n18829), .Y(n19986) );
  xor2_1 U19775 ( .A(n19987), .B(n18682), .X(n18829) );
  nand2_1 U19776 ( .A(n13031), .B(n19988), .Y(n19987) );
  xnor2_1 U19777 ( .A(n19989), .B(n11751), .Y(n18826) );
  o22ai_1 U19778 ( .A1(n19990), .A2(n16314), .B1(n19991), .B2(n17000), .Y(
        n19989) );
  inv_1 U19779 ( .A(n23884), .Y(n17000) );
  nor2_1 U19780 ( .A(n11763), .B(n19975), .Y(n19991) );
  inv_1 U19781 ( .A(n11763), .Y(n16314) );
  xor2_1 U19782 ( .A(n19992), .B(n19993), .X(n11763) );
  xor2_1 U19783 ( .A(n19994), .B(n18466), .X(n19993) );
  inv_1 U19784 ( .A(n17765), .Y(n18466) );
  xor2_1 U19785 ( .A(n15953), .B(n12380), .X(n19992) );
  inv_1 U19786 ( .A(n19975), .Y(n19990) );
  o22ai_1 U19787 ( .A1(n11631), .A2(n19181), .B1(n12446), .B2(n19995), .Y(
        n19975) );
  nor2_1 U19788 ( .A(n19996), .B(n16307), .Y(n19995) );
  inv_1 U19789 ( .A(n19996), .Y(n19181) );
  a21oi_1 U19790 ( .A1(n19177), .A2(n12445), .B1(n19179), .Y(n19996) );
  a211oi_1 U19791 ( .A1(n19170), .A2(n17003), .B1(n19997), .C1(n16872), .Y(
        n19179) );
  a21oi_1 U19792 ( .A1(n16277), .A2(n19998), .B1(n1519), .Y(n19997) );
  o211ai_1 U19793 ( .A1(n17003), .A2(n19170), .B1(n19999), .C1(n16872), .Y(
        n19177) );
  xor2_1 U19794 ( .A(n20000), .B(n20001), .X(n16872) );
  xor2_1 U19795 ( .A(n20002), .B(n11294), .X(n20001) );
  inv_1 U19796 ( .A(n18034), .Y(n11294) );
  xor2_1 U19797 ( .A(n13010), .B(n20003), .X(n20000) );
  xor2_1 U19798 ( .A(n23950), .B(n12299), .X(n20003) );
  nand3_1 U19799 ( .A(n20004), .B(n20005), .C(n20006), .Y(n13010) );
  o21ai_0 U19800 ( .A1(n19865), .A2(n19864), .B1(n24027), .Y(n20006) );
  o211ai_1 U19801 ( .A1(n24028), .A2(n20007), .B1(n12416), .C1(n19318), .Y(
        n20004) );
  o21ai_0 U19802 ( .A1(n19998), .A2(n16277), .B1(n1519), .Y(n19999) );
  inv_1 U19803 ( .A(n17003), .Y(n16277) );
  inv_1 U19804 ( .A(n19998), .Y(n19170) );
  xor2_1 U19805 ( .A(n20008), .B(n16222), .X(n19998) );
  o22ai_1 U19806 ( .A1(n20009), .A2(n18111), .B1(n12515), .B2(n20010), .Y(
        n20008) );
  nor2_1 U19807 ( .A(n18110), .B(n18870), .Y(n20010) );
  inv_1 U19808 ( .A(n18110), .Y(n18111) );
  xnor2_1 U19809 ( .A(n17992), .B(n16882), .Y(n18110) );
  inv_1 U19810 ( .A(n12879), .Y(n16882) );
  xnor2_1 U19811 ( .A(n20011), .B(n20012), .Y(n12879) );
  xor2_1 U19812 ( .A(n18305), .B(n12320), .X(n20011) );
  nand4_1 U19813 ( .A(n12359), .B(n20013), .C(n20014), .D(n20015), .Y(n17992)
         );
  a211oi_1 U19814 ( .A1(n19318), .A2(n20016), .B1(n20017), .C1(n20018), .Y(
        n20015) );
  inv_1 U19815 ( .A(n19858), .Y(n20018) );
  a21oi_1 U19816 ( .A1(n20019), .A2(n24027), .B1(n12339), .Y(n19858) );
  o21ai_0 U19817 ( .A1(n12416), .A2(n20020), .B1(n20005), .Y(n20019) );
  mux2_1 U19818 ( .A0(n12419), .A1(n12338), .S(n12407), .X(n20017) );
  nor2_1 U19819 ( .A(n20021), .B(n10610), .Y(n12338) );
  nor2_1 U19820 ( .A(n12370), .B(n24029), .Y(n12419) );
  nor2_1 U19821 ( .A(n20020), .B(n24027), .Y(n19318) );
  nand3_1 U19822 ( .A(n12387), .B(n10610), .C(n19317), .Y(n20014) );
  nand2_1 U19823 ( .A(n19864), .B(n24030), .Y(n12359) );
  inv_1 U19824 ( .A(n18870), .Y(n20009) );
  o21ai_0 U19825 ( .A1(n12890), .A2(n12894), .B1(n20022), .Y(n18870) );
  xor2_1 U19826 ( .A(n24045), .B(n20023), .X(n20022) );
  nor2_1 U19827 ( .A(n19156), .B(n19157), .Y(n20023) );
  a21oi_1 U19828 ( .A1(n10623), .A2(n16637), .B1(n20024), .Y(n19157) );
  xor2_1 U19829 ( .A(n23903), .B(n20025), .X(n20024) );
  or2_0 U19830 ( .A(n18892), .B(n18891), .X(n20025) );
  nor2_1 U19831 ( .A(n10623), .B(n16637), .Y(n18891) );
  inv_1 U19832 ( .A(n18893), .Y(n18892) );
  o21ai_0 U19833 ( .A1(n18905), .A2(n18908), .B1(n18907), .Y(n18893) );
  nand2_1 U19834 ( .A(n16625), .B(n10644), .Y(n18907) );
  xor2_1 U19835 ( .A(n17611), .B(n20026), .X(n18908) );
  nor2_1 U19836 ( .A(n16625), .B(n10644), .Y(n20026) );
  inv_1 U19837 ( .A(n12907), .Y(n16625) );
  xnor2_1 U19838 ( .A(n20027), .B(n17598), .Y(n12907) );
  o211ai_1 U19839 ( .A1(n14707), .A2(n14696), .B1(n20028), .C1(n20029), .Y(
        n17598) );
  a222oi_1 U19840 ( .A1(n19142), .A2(n20030), .B1(n14682), .B2(n20031), .C1(
        n14596), .C2(n20032), .Y(n20029) );
  o22ai_1 U19841 ( .A1(n24017), .A2(n20030), .B1(n24047), .B2(n14675), .Y(
        n20032) );
  nand2_1 U19842 ( .A(n14695), .B(n14625), .Y(n20031) );
  inv_1 U19843 ( .A(n14665), .Y(n14682) );
  nand2_1 U19844 ( .A(n24039), .B(n20033), .Y(n14665) );
  xnor2_1 U19845 ( .A(n20034), .B(n20035), .Y(n20027) );
  nand2_1 U19846 ( .A(n20036), .B(n20037), .Y(n20034) );
  inv_1 U19847 ( .A(n20038), .Y(n20037) );
  a21oi_1 U19848 ( .A1(n20039), .A2(n16516), .B1(n20040), .Y(n18905) );
  a21oi_1 U19849 ( .A1(n17761), .A2(n19147), .B1(n17356), .Y(n20040) );
  inv_1 U19850 ( .A(n23702), .Y(n17356) );
  inv_1 U19851 ( .A(n16516), .Y(n17761) );
  xor2_1 U19852 ( .A(n20041), .B(n20042), .X(n16516) );
  xor2_1 U19853 ( .A(n23958), .B(n23948), .X(n20042) );
  xnor2_1 U19854 ( .A(n20043), .B(n17152), .Y(n20041) );
  inv_1 U19855 ( .A(n19147), .Y(n20039) );
  xor2_1 U19856 ( .A(n20044), .B(n18724), .X(n19147) );
  inv_1 U19857 ( .A(n17458), .Y(n18724) );
  o221ai_1 U19858 ( .A1(n20045), .A2(n10616), .B1(n16140), .B2(n20046), .C1(
        n20047), .Y(n17458) );
  a21oi_1 U19859 ( .A1(n23962), .A2(n20048), .B1(n20049), .Y(n20047) );
  mux2i_1 U19860 ( .A0(n16189), .A1(n20050), .S(n23960), .Y(n20049) );
  nand2_1 U19861 ( .A(n20051), .B(n16155), .Y(n20050) );
  o22ai_1 U19862 ( .A1(n23961), .A2(n20052), .B1(n16100), .B2(n16144), .Y(
        n20048) );
  o22ai_1 U19863 ( .A1(n16542), .A2(n20053), .B1(n2116), .B2(n20054), .Y(
        n20044) );
  nor2_1 U19864 ( .A(n19127), .B(n16906), .Y(n20054) );
  inv_1 U19865 ( .A(n16542), .Y(n16906) );
  inv_1 U19866 ( .A(n19127), .Y(n20053) );
  xor2_1 U19867 ( .A(n20055), .B(n12297), .X(n19127) );
  o22ai_1 U19868 ( .A1(n16550), .A2(n18925), .B1(n23676), .B2(n20056), .Y(
        n20055) );
  and2_0 U19869 ( .A(n18925), .B(n16550), .X(n20056) );
  mux2i_1 U19870 ( .A0(n19121), .A1(n20057), .S(n19507), .Y(n18925) );
  a21oi_1 U19871 ( .A1(n19123), .A2(n19124), .B1(n20058), .Y(n20057) );
  inv_1 U19872 ( .A(n19122), .Y(n20058) );
  and3_1 U19873 ( .A(n19123), .B(n19122), .C(n19124), .X(n19121) );
  xnor2_1 U19874 ( .A(n13410), .B(n20059), .Y(n19124) );
  a21oi_1 U19875 ( .A1(n19108), .A2(n19110), .B1(n19111), .Y(n20059) );
  xor2_1 U19876 ( .A(n19009), .B(n20060), .X(n19111) );
  nor2_1 U19877 ( .A(n23826), .B(n16916), .Y(n20060) );
  nand2_1 U19878 ( .A(n23826), .B(n16916), .Y(n19110) );
  xor2_1 U19879 ( .A(n20061), .B(n23958), .X(n16916) );
  nand2_1 U19880 ( .A(n20062), .B(n20063), .Y(n20061) );
  o21ai_0 U19881 ( .A1(n19106), .A2(n16921), .B1(n19105), .Y(n19108) );
  nand2_1 U19882 ( .A(n20064), .B(n11388), .Y(n19105) );
  inv_1 U19883 ( .A(n16583), .Y(n16921) );
  xor2_1 U19884 ( .A(n20065), .B(n20066), .X(n16583) );
  xor2_1 U19885 ( .A(n23981), .B(n12393), .X(n20066) );
  xor2_1 U19886 ( .A(n20067), .B(n16914), .X(n20065) );
  inv_1 U19887 ( .A(n16493), .Y(n16914) );
  o21ai_0 U19888 ( .A1(n20068), .A2(n20069), .B1(n13392), .Y(n16493) );
  mux2i_1 U19889 ( .A0(n13398), .A1(n23982), .S(n24013), .Y(n20069) );
  nor2_1 U19890 ( .A(n11388), .B(n20064), .Y(n19106) );
  a22oi_1 U19891 ( .A1(n19097), .A2(n16507), .B1(n20070), .B2(n12442), .Y(
        n20064) );
  or2_0 U19892 ( .A(n16507), .B(n19097), .X(n20070) );
  inv_1 U19893 ( .A(n17777), .Y(n16507) );
  xor2_1 U19894 ( .A(n20071), .B(n20072), .X(n17777) );
  xor2_1 U19895 ( .A(n11168), .B(n20073), .X(n20072) );
  xor2_1 U19896 ( .A(n10606), .B(n12394), .X(n20071) );
  o22ai_1 U19897 ( .A1(n16482), .A2(n18949), .B1(n20074), .B2(n12711), .Y(
        n19097) );
  inv_1 U19898 ( .A(n23857), .Y(n12711) );
  and2_0 U19899 ( .A(n18949), .B(n16482), .X(n20074) );
  o22ai_1 U19900 ( .A1(n20075), .A2(n16925), .B1(n20076), .B2(n12718), .Y(
        n18949) );
  inv_1 U19901 ( .A(n23767), .Y(n12718) );
  nor2_1 U19902 ( .A(n12705), .B(n18952), .Y(n20076) );
  inv_1 U19903 ( .A(n12705), .Y(n16925) );
  xor2_1 U19904 ( .A(n20077), .B(n20078), .X(n12705) );
  a21oi_1 U19905 ( .A1(n20079), .A2(n18040), .B1(n20080), .Y(n20078) );
  a21oi_1 U19906 ( .A1(n23985), .A2(n15990), .B1(n20081), .Y(n20079) );
  inv_1 U19907 ( .A(n20082), .Y(n20081) );
  inv_1 U19908 ( .A(n18952), .Y(n20075) );
  o22ai_1 U19909 ( .A1(n12715), .A2(n19095), .B1(n23864), .B2(n20083), .Y(
        n18952) );
  and2_0 U19910 ( .A(n19095), .B(n12715), .X(n20083) );
  o22ai_1 U19911 ( .A1(n11130), .A2(n20084), .B1(n23865), .B2(n20085), .Y(
        n19095) );
  nor2_1 U19912 ( .A(n19085), .B(n16933), .Y(n20085) );
  inv_1 U19913 ( .A(n11130), .Y(n16933) );
  inv_1 U19914 ( .A(n19085), .Y(n20084) );
  xor2_1 U19915 ( .A(n20086), .B(n18021), .X(n19085) );
  inv_1 U19916 ( .A(n18358), .Y(n18021) );
  nand3_1 U19917 ( .A(n20087), .B(n20088), .C(n20089), .Y(n18358) );
  a221oi_1 U19918 ( .A1(n23977), .A2(n19411), .B1(n16071), .B2(n20090), .C1(
        n20091), .Y(n20089) );
  inv_1 U19919 ( .A(n19952), .Y(n20091) );
  nand3_1 U19920 ( .A(n16134), .B(n16163), .C(n23974), .Y(n19952) );
  o21ai_0 U19921 ( .A1(n23975), .A2(n19415), .B1(n20092), .Y(n20090) );
  a22oi_1 U19922 ( .A1(n18844), .A2(n19414), .B1(n18843), .B2(n20093), .Y(
        n20087) );
  o21ai_0 U19923 ( .A1(n19073), .A2(n12725), .B1(n19071), .Y(n20086) );
  nand2_1 U19924 ( .A(n20748), .B(n20094), .Y(n19071) );
  xor2_1 U19925 ( .A(n20095), .B(n20096), .X(n12725) );
  mux2i_1 U19926 ( .A0(n20097), .A1(n20098), .S(n12401), .Y(n20096) );
  nand2_1 U19927 ( .A(n16995), .B(n20099), .Y(n20098) );
  nand2_1 U19928 ( .A(n11751), .B(n20100), .Y(n20097) );
  nor2_1 U19929 ( .A(n20094), .B(n20748), .Y(n19073) );
  xor2_1 U19930 ( .A(n18034), .B(n20101), .X(n20094) );
  o21ai_0 U19931 ( .A1(n19062), .A2(n19065), .B1(n19063), .Y(n20101) );
  xnor2_1 U19932 ( .A(n12817), .B(n20102), .Y(n19063) );
  nor2_1 U19933 ( .A(n23709), .B(n11136), .Y(n20102) );
  nor2_1 U19934 ( .A(n11118), .B(n16938), .Y(n19065) );
  inv_1 U19935 ( .A(n11136), .Y(n16938) );
  xor2_1 U19936 ( .A(n20103), .B(n20104), .X(n11136) );
  xor2_1 U19937 ( .A(n20105), .B(n18136), .X(n20103) );
  inv_1 U19938 ( .A(n23709), .Y(n11118) );
  a21oi_1 U19939 ( .A1(n16940), .A2(n23867), .B1(n20106), .Y(n19062) );
  xor2_1 U19940 ( .A(n12984), .B(n20107), .X(n20106) );
  o21ai_0 U19941 ( .A1(n23867), .A2(n16940), .B1(n18975), .Y(n20107) );
  xor2_1 U19942 ( .A(n20108), .B(n12297), .X(n18975) );
  o22ai_1 U19943 ( .A1(n20109), .A2(n19059), .B1(n2122), .B2(n20110), .Y(
        n20108) );
  nor2_1 U19944 ( .A(n12731), .B(n19058), .Y(n20110) );
  inv_1 U19945 ( .A(n16674), .Y(n12731) );
  xnor2_1 U19946 ( .A(n16674), .B(n17737), .Y(n19059) );
  xor2_1 U19947 ( .A(n20111), .B(n20112), .X(n16674) );
  xor2_1 U19948 ( .A(n24022), .B(n12305), .X(n20112) );
  inv_1 U19949 ( .A(n19058), .Y(n20109) );
  o21ai_0 U19950 ( .A1(n16414), .A2(n20113), .B1(n20114), .Y(n19058) );
  o21ai_0 U19951 ( .A1(n19051), .A2(n16415), .B1(n23869), .Y(n20114) );
  inv_1 U19952 ( .A(n20113), .Y(n19051) );
  o21ai_0 U19953 ( .A1(n23863), .A2(n11120), .B1(n20115), .Y(n20113) );
  xor2_1 U19954 ( .A(n11742), .B(n20116), .X(n20115) );
  a21oi_1 U19955 ( .A1(n23863), .A2(n11120), .B1(n19044), .Y(n20116) );
  o22ai_1 U19956 ( .A1(n19006), .A2(n16391), .B1(n23882), .B2(n20117), .Y(
        n19044) );
  nor2_1 U19957 ( .A(n16947), .B(n20118), .Y(n20117) );
  inv_1 U19958 ( .A(n16391), .Y(n16947) );
  xor2_1 U19959 ( .A(n20119), .B(n20120), .X(n16391) );
  xor2_1 U19960 ( .A(n15880), .B(n24011), .X(n20119) );
  inv_1 U19961 ( .A(n20118), .Y(n19006) );
  nand2_1 U19962 ( .A(n18738), .B(n11531), .Y(n20118) );
  xnor2_1 U19963 ( .A(n20121), .B(n20122), .Y(n11531) );
  a21oi_1 U19964 ( .A1(n12331), .A2(n24022), .B1(n20123), .Y(n20122) );
  nor2_1 U19965 ( .A(n17966), .B(n20124), .Y(n18738) );
  nand3_1 U19966 ( .A(n15880), .B(n10609), .C(n12333), .Y(n17966) );
  inv_1 U19967 ( .A(n17860), .Y(n11742) );
  inv_1 U19968 ( .A(n17793), .Y(n11120) );
  xnor2_1 U19969 ( .A(n20125), .B(n20126), .Y(n17793) );
  nor2_1 U19970 ( .A(n20127), .B(n20128), .Y(n20126) );
  xor2_1 U19971 ( .A(n16222), .B(n20129), .X(n20128) );
  inv_1 U19972 ( .A(n16832), .Y(n16222) );
  o21ai_0 U19973 ( .A1(n20130), .A2(n20131), .B1(n19814), .Y(n16832) );
  inv_1 U19974 ( .A(n20132), .Y(n20127) );
  inv_1 U19975 ( .A(n16415), .Y(n16414) );
  xor2_1 U19976 ( .A(n20133), .B(n20134), .X(n16415) );
  xor2_1 U19977 ( .A(n16627), .B(n20135), .X(n20134) );
  o221ai_1 U19978 ( .A1(n20045), .A2(n20046), .B1(n23962), .B2(n20136), .C1(
        n20137), .Y(n16627) );
  a211oi_1 U19979 ( .A1(n16137), .A2(n23963), .B1(n16062), .C1(n16037), .Y(
        n20137) );
  inv_1 U19980 ( .A(n16167), .Y(n16037) );
  nand2_1 U19981 ( .A(n20051), .B(n16100), .Y(n16167) );
  inv_1 U19982 ( .A(n16166), .Y(n16062) );
  nand2_1 U19983 ( .A(n16172), .B(n16162), .Y(n16166) );
  mux2i_1 U19984 ( .A0(n16162), .A1(n16087), .S(n16088), .Y(n20136) );
  mux2i_1 U19985 ( .A0(n16168), .A1(n16100), .S(n23962), .Y(n20045) );
  o211ai_1 U19986 ( .A1(n12333), .A2(n13401), .B1(n20138), .C1(n20139), .Y(
        n20133) );
  o21ai_0 U19987 ( .A1(n13307), .A2(n15920), .B1(n18463), .Y(n20138) );
  xor2_1 U19988 ( .A(n20140), .B(n20141), .X(n16940) );
  o221ai_1 U19989 ( .A1(n23983), .A2(n13404), .B1(n24013), .B2(n13403), .C1(
        n20142), .Y(n18034) );
  a211oi_1 U19990 ( .A1(n20068), .A2(n18672), .B1(n13350), .C1(n13308), .Y(
        n20142) );
  nor2_1 U19991 ( .A(n13392), .B(n13378), .Y(n13308) );
  nor2_1 U19992 ( .A(n13379), .B(n13382), .Y(n13350) );
  xor2_1 U19993 ( .A(n20143), .B(n20144), .X(n11130) );
  nor2_1 U19994 ( .A(n20145), .B(n20146), .Y(n20144) );
  xor2_1 U19995 ( .A(n20147), .B(n20148), .X(n12715) );
  xnor2_1 U19996 ( .A(n20149), .B(n20150), .Y(n16482) );
  xor2_1 U19997 ( .A(n16510), .B(n23987), .X(n20149) );
  inv_1 U19998 ( .A(n12582), .Y(n11388) );
  nand2_1 U19999 ( .A(n20151), .B(n17326), .Y(n19122) );
  xor2_1 U20000 ( .A(n17525), .B(n16912), .X(n20151) );
  inv_1 U20001 ( .A(n18066), .Y(n17525) );
  xnor2_1 U20002 ( .A(n11413), .B(n20152), .Y(n19123) );
  nor2_1 U20003 ( .A(n16912), .B(n17326), .Y(n20152) );
  inv_1 U20004 ( .A(n12581), .Y(n17326) );
  xor2_1 U20005 ( .A(n20153), .B(n20154), .X(n16912) );
  nand2_1 U20006 ( .A(n20155), .B(n20156), .Y(n20153) );
  xor2_1 U20007 ( .A(n20157), .B(n20158), .X(n16550) );
  a21oi_1 U20008 ( .A1(n20159), .A2(n17479), .B1(n20160), .Y(n20158) );
  a21oi_1 U20009 ( .A1(n16524), .A2(n10606), .B1(n20161), .Y(n20159) );
  xor2_1 U20010 ( .A(n20162), .B(n20163), .X(n16542) );
  xor2_1 U20011 ( .A(n15902), .B(n12302), .X(n20162) );
  xor2_1 U20012 ( .A(n20164), .B(n20165), .X(n16637) );
  o211ai_1 U20013 ( .A1(n12299), .A2(n17310), .B1(n20166), .C1(n20167), .Y(
        n20164) );
  o21ai_0 U20014 ( .A1(n12629), .A2(n15955), .B1(n12319), .Y(n20166) );
  nor2_1 U20015 ( .A(n16894), .B(n8), .Y(n19156) );
  inv_1 U20016 ( .A(n12890), .Y(n16894) );
  inv_1 U20017 ( .A(n8), .Y(n12894) );
  xor2_1 U20018 ( .A(n20168), .B(n20169), .X(n12890) );
  xor2_1 U20019 ( .A(n20170), .B(n11205), .X(n20169) );
  inv_1 U20020 ( .A(n11346), .Y(n11205) );
  xor2_1 U20021 ( .A(n20171), .B(n20172), .X(n17003) );
  xor2_1 U20022 ( .A(n23953), .B(n23938), .X(n20172) );
  xnor2_1 U20023 ( .A(n20173), .B(n17746), .Y(n20171) );
  inv_1 U20024 ( .A(n16307), .Y(n11631) );
  xor2_1 U20025 ( .A(n20174), .B(n23951), .X(n16307) );
  o21ai_0 U20026 ( .A1(n20175), .A2(n16015), .B1(n20176), .Y(n20174) );
  nor2_1 U20027 ( .A(n19988), .B(n13031), .Y(n18828) );
  inv_1 U20028 ( .A(n16863), .Y(n13031) );
  o21ai_0 U20029 ( .A1(n16013), .A2(n20177), .B1(n20178), .Y(n16863) );
  mux2i_1 U20030 ( .A0(n20179), .A1(n20180), .S(n12380), .Y(n20178) );
  inv_1 U20031 ( .A(n19984), .Y(n20180) );
  nor2_1 U20032 ( .A(n23938), .B(n20181), .Y(n20179) );
  xor2_1 U20033 ( .A(n10826), .B(n20181), .X(n20177) );
  inv_1 U20034 ( .A(n12522), .Y(n19988) );
  nand2_1 U20035 ( .A(n18767), .B(n20182), .Y(n19976) );
  inv_1 U20036 ( .A(n18768), .Y(n20182) );
  nor2_1 U20037 ( .A(n16229), .B(n818), .Y(n18768) );
  xnor2_1 U20038 ( .A(n10879), .B(n20183), .Y(n18767) );
  and2_0 U20039 ( .A(n16229), .B(n818), .X(n20183) );
  inv_1 U20040 ( .A(n16226), .Y(n16229) );
  mux2i_1 U20041 ( .A0(n20184), .A1(n20185), .S(n18682), .Y(n16226) );
  inv_1 U20042 ( .A(n17591), .Y(n18682) );
  o211ai_1 U20043 ( .A1(n12403), .A2(n12396), .B1(n20186), .C1(n20187), .Y(
        n17591) );
  xnor2_1 U20044 ( .A(n18763), .B(n20188), .Y(n20185) );
  xor2_1 U20045 ( .A(n18763), .B(n18764), .X(n20184) );
  xnor2_1 U20046 ( .A(n20189), .B(n17697), .Y(n18763) );
  inv_1 U20047 ( .A(n17988), .Y(n17697) );
  o21ai_0 U20048 ( .A1(n24032), .A2(n12356), .B1(n20190), .Y(n17988) );
  mux2i_1 U20049 ( .A0(n12390), .A1(n19875), .S(n19529), .Y(n20190) );
  nand2_1 U20050 ( .A(n12384), .B(n24026), .Y(n12356) );
  o221ai_1 U20051 ( .A1(n10607), .A2(n19984), .B1(n20191), .B2(n19982), .C1(
        n19985), .Y(n20189) );
  o21ai_0 U20052 ( .A1(n20181), .A2(n16013), .B1(n10826), .Y(n19985) );
  xnor2_1 U20053 ( .A(n16275), .B(n20192), .Y(n19982) );
  nor2_1 U20054 ( .A(n12380), .B(n10607), .Y(n20192) );
  nand4_1 U20055 ( .A(n20193), .B(n18873), .C(n18874), .D(n12385), .Y(n16275)
         );
  inv_1 U20056 ( .A(n19684), .Y(n18873) );
  mux2i_1 U20057 ( .A0(n12222), .A1(n12422), .S(n24025), .Y(n20193) );
  inv_1 U20058 ( .A(n19981), .Y(n20191) );
  nand2_1 U20059 ( .A(n20181), .B(n16013), .Y(n19984) );
  xor2_1 U20060 ( .A(n20194), .B(n11346), .X(n20181) );
  nor4_1 U20061 ( .A(n20195), .B(n13743), .C(n13838), .D(n13725), .Y(n11346)
         );
  and2_0 U20062 ( .A(n13921), .B(n13927), .X(n13838) );
  nor2_1 U20063 ( .A(n19970), .B(n13947), .Y(n13743) );
  and2_0 U20064 ( .A(n13926), .B(n23999), .X(n20195) );
  o22ai_1 U20065 ( .A1(n15953), .A2(n19994), .B1(n20196), .B2(n10826), .Y(
        n20194) );
  and2_0 U20066 ( .A(n19994), .B(n15953), .X(n20196) );
  nand2_1 U20067 ( .A(n20176), .B(n20197), .Y(n19994) );
  o21ai_0 U20068 ( .A1(n20175), .A2(n16015), .B1(n23951), .Y(n20197) );
  nand2_1 U20069 ( .A(n20175), .B(n16015), .Y(n20176) );
  xnor2_1 U20070 ( .A(n20198), .B(n17152), .Y(n20175) );
  o22ai_1 U20071 ( .A1(n12299), .A2(n20002), .B1(n23950), .B2(n20199), .Y(
        n20198) );
  nor2_1 U20072 ( .A(n15955), .B(n20200), .Y(n20199) );
  inv_1 U20073 ( .A(n20200), .Y(n20002) );
  o22ai_1 U20074 ( .A1(n16013), .A2(n20173), .B1(n20201), .B2(n16611), .Y(
        n20200) );
  and2_0 U20075 ( .A(n20173), .B(n16013), .X(n20201) );
  o22ai_1 U20076 ( .A1(n12320), .A2(n20012), .B1(n20202), .B2(n18305), .Y(
        n20173) );
  and2_0 U20077 ( .A(n20012), .B(n12320), .X(n20202) );
  mux2i_1 U20078 ( .A0(n20203), .A1(n20204), .S(n10946), .Y(n20012) );
  a21oi_1 U20079 ( .A1(n20205), .A2(n20206), .B1(n20207), .Y(n20204) );
  inv_1 U20080 ( .A(n20208), .Y(n20207) );
  inv_1 U20081 ( .A(n20168), .Y(n20205) );
  nor2_1 U20082 ( .A(n20168), .B(n20170), .Y(n20203) );
  nand2_1 U20083 ( .A(n20206), .B(n20208), .Y(n20170) );
  nand2_1 U20084 ( .A(n12302), .B(n20209), .Y(n20208) );
  xor2_1 U20085 ( .A(n20210), .B(n11520), .X(n20206) );
  nand2_1 U20086 ( .A(n23951), .B(n15931), .Y(n20210) );
  o221ai_1 U20087 ( .A1(n20211), .A2(n15955), .B1(n12319), .B2(n20212), .C1(
        n20167), .Y(n20168) );
  nand3_1 U20088 ( .A(n17310), .B(n16524), .C(n12299), .Y(n20167) );
  inv_1 U20089 ( .A(n12629), .Y(n17310) );
  a21oi_1 U20090 ( .A1(n12629), .A2(n15955), .B1(n20213), .Y(n20212) );
  a21oi_1 U20091 ( .A1(n12319), .A2(n12629), .B1(n20213), .Y(n20211) );
  inv_1 U20092 ( .A(n20165), .Y(n20213) );
  o21ai_0 U20093 ( .A1(n20038), .A2(n20035), .B1(n20036), .Y(n20165) );
  xor2_1 U20094 ( .A(n20214), .B(n14685), .X(n20036) );
  nand2_1 U20095 ( .A(n23959), .B(n23953), .Y(n20214) );
  o22ai_1 U20096 ( .A1(n20043), .A2(n18305), .B1(n20215), .B2(n18413), .Y(
        n20035) );
  and2_0 U20097 ( .A(n20043), .B(n18305), .X(n20215) );
  o22ai_1 U20098 ( .A1(n15931), .A2(n20216), .B1(n12393), .B2(n20217), .Y(
        n20043) );
  nor2_1 U20099 ( .A(n20163), .B(n12302), .Y(n20217) );
  inv_1 U20100 ( .A(n20163), .Y(n20216) );
  a22oi_1 U20101 ( .A1(n20218), .A2(n20160), .B1(n20219), .B2(n17479), .Y(
        n20163) );
  o22ai_1 U20102 ( .A1(n20157), .A2(n20161), .B1(n12319), .B2(n1965), .Y(
        n20219) );
  and2_0 U20103 ( .A(n20161), .B(n18086), .X(n20160) );
  inv_1 U20104 ( .A(n17479), .Y(n18086) );
  nor3_1 U20105 ( .A(n18443), .B(n13939), .C(n20220), .Y(n17479) );
  o22ai_1 U20106 ( .A1(n18445), .A2(n20221), .B1(n1678), .B2(n24009), .Y(
        n20220) );
  inv_1 U20107 ( .A(n24008), .Y(n20221) );
  nor2_1 U20108 ( .A(n10606), .B(n16524), .Y(n20161) );
  inv_1 U20109 ( .A(n20157), .Y(n20218) );
  nand2_1 U20110 ( .A(n20155), .B(n20222), .Y(n20157) );
  xor2_1 U20111 ( .A(n13410), .B(n20223), .X(n20222) );
  nand2_1 U20112 ( .A(n20154), .B(n20156), .Y(n20223) );
  nand2_1 U20113 ( .A(n16545), .B(n16510), .Y(n20156) );
  a21oi_1 U20114 ( .A1(n20062), .A2(n23958), .B1(n20224), .Y(n20154) );
  inv_1 U20115 ( .A(n20063), .Y(n20224) );
  o211ai_1 U20116 ( .A1(n12393), .A2(n20225), .B1(n20226), .C1(n15990), .Y(
        n20063) );
  o21ai_0 U20117 ( .A1(n20067), .A2(n15902), .B1(n15999), .Y(n20226) );
  o211ai_1 U20118 ( .A1(n20067), .A2(n15902), .B1(n20227), .C1(n12392), .Y(
        n20062) );
  o21ai_0 U20119 ( .A1(n20225), .A2(n12393), .B1(n23981), .Y(n20227) );
  inv_1 U20120 ( .A(n20067), .Y(n20225) );
  o22ai_1 U20121 ( .A1(n20228), .A2(n15992), .B1(n20229), .B2(n10606), .Y(
        n20067) );
  nor2_1 U20122 ( .A(n12394), .B(n20073), .Y(n20229) );
  inv_1 U20123 ( .A(n20073), .Y(n20228) );
  o22ai_1 U20124 ( .A1(n16510), .A2(n20150), .B1(n20230), .B2(n16453), .Y(
        n20073) );
  and2_0 U20125 ( .A(n20150), .B(n16510), .X(n20230) );
  o32ai_1 U20126 ( .A1(n18262), .A2(n12392), .A3(n16464), .B1(n20231), .B2(
        n20077), .Y(n20150) );
  xor2_1 U20127 ( .A(n12686), .B(n20232), .X(n20077) );
  mux2i_1 U20128 ( .A0(n20233), .A1(n20234), .S(n20235), .Y(n20232) );
  inv_1 U20129 ( .A(n17133), .Y(n20235) );
  o221ai_1 U20130 ( .A1(n13384), .A2(n13367), .B1(n24003), .B2(n19560), .C1(
        n13369), .Y(n17133) );
  o22ai_1 U20131 ( .A1(n20236), .A2(n15999), .B1(n12388), .B2(n20237), .Y(
        n20234) );
  nor2_1 U20132 ( .A(n20148), .B(n23981), .Y(n20237) );
  inv_1 U20133 ( .A(n20148), .Y(n20236) );
  nor2_1 U20134 ( .A(n20148), .B(n20147), .Y(n20233) );
  xor2_1 U20135 ( .A(n15970), .B(n15999), .X(n20147) );
  nor2_1 U20136 ( .A(n20146), .B(n20238), .Y(n20148) );
  xor2_1 U20137 ( .A(n11413), .B(n20239), .X(n20238) );
  nor2_1 U20138 ( .A(n20145), .B(n20143), .Y(n20239) );
  nand2_1 U20139 ( .A(n20240), .B(n20241), .Y(n20143) );
  nand3_1 U20140 ( .A(n11489), .B(n18463), .C(n20100), .Y(n20241) );
  xor2_1 U20141 ( .A(n16995), .B(n23987), .X(n20100) );
  mux2i_1 U20142 ( .A0(n20242), .A1(n20243), .S(n16995), .Y(n20240) );
  a221oi_1 U20143 ( .A1(n12407), .A2(n20244), .B1(n20016), .B2(n19317), .C1(
        n19861), .Y(n16995) );
  nor3_1 U20144 ( .A(n12407), .B(n24028), .C(n12374), .Y(n19861) );
  nor2_1 U20145 ( .A(n12407), .B(n24024), .Y(n19317) );
  or3_1 U20146 ( .A(n12339), .B(n12267), .C(n12336), .X(n20244) );
  nor3_1 U20147 ( .A(n20020), .B(n24029), .C(n12428), .Y(n12336) );
  inv_1 U20148 ( .A(n24024), .Y(n20020) );
  inv_1 U20149 ( .A(n20245), .Y(n12267) );
  nor2_1 U20150 ( .A(n20005), .B(n24029), .Y(n12339) );
  o22ai_1 U20151 ( .A1(n20099), .A2(n18463), .B1(n20246), .B2(n20095), .Y(
        n20243) );
  inv_1 U20152 ( .A(n20247), .Y(n20246) );
  xor2_1 U20153 ( .A(n11489), .B(n23987), .X(n20099) );
  nor2_1 U20154 ( .A(n20095), .B(n20247), .Y(n20242) );
  nand2_1 U20155 ( .A(n23987), .B(n18463), .Y(n20247) );
  mux2i_1 U20156 ( .A0(n20248), .A1(n20249), .S(n17915), .Y(n20095) );
  inv_1 U20157 ( .A(n19817), .Y(n17915) );
  o221ai_1 U20158 ( .A1(n14695), .A2(n14687), .B1(n24038), .B2(n14663), .C1(
        n20250), .Y(n19817) );
  a21oi_1 U20159 ( .A1(n19671), .A2(n20251), .B1(n19142), .Y(n20250) );
  nor2_1 U20160 ( .A(n14702), .B(n14676), .Y(n19142) );
  nand2_1 U20161 ( .A(n24046), .B(n14707), .Y(n20251) );
  nand3_1 U20162 ( .A(n20252), .B(n14676), .C(n24046), .Y(n14695) );
  a21oi_1 U20163 ( .A1(n20104), .A2(n20253), .B1(n20254), .Y(n20249) );
  inv_1 U20164 ( .A(n20255), .Y(n20254) );
  inv_1 U20165 ( .A(n20256), .Y(n20104) );
  nor2_1 U20166 ( .A(n20256), .B(n20105), .Y(n20248) );
  nand2_1 U20167 ( .A(n20253), .B(n20255), .Y(n20105) );
  nand2_1 U20168 ( .A(n23993), .B(n18262), .Y(n20255) );
  xor2_1 U20169 ( .A(n12530), .B(n20257), .X(n20253) );
  nor2_1 U20170 ( .A(n23993), .B(n18262), .Y(n20257) );
  inv_1 U20171 ( .A(n16535), .Y(n12530) );
  nand4_1 U20172 ( .A(n12409), .B(n12334), .C(n12404), .D(n18874), .Y(n16535)
         );
  nand2_1 U20173 ( .A(n12421), .B(n20258), .Y(n18874) );
  inv_1 U20174 ( .A(n12396), .Y(n12421) );
  mux2i_1 U20175 ( .A0(n20259), .A1(n20260), .S(n18588), .Y(n20256) );
  inv_1 U20176 ( .A(n11525), .Y(n18588) );
  mux2i_1 U20177 ( .A0(n14661), .A1(n14683), .S(n24042), .Y(n11525) );
  nand2_1 U20178 ( .A(n20261), .B(n20141), .Y(n20260) );
  xor2_1 U20179 ( .A(n24011), .B(n12388), .X(n20141) );
  o22ai_1 U20180 ( .A1(n10608), .A2(n20140), .B1(n20262), .B2(n15970), .Y(
        n20259) );
  nor2_1 U20181 ( .A(n20261), .B(n24011), .Y(n20262) );
  inv_1 U20182 ( .A(n20140), .Y(n20261) );
  o22ai_1 U20183 ( .A1(n12305), .A2(n20263), .B1(n24022), .B2(n20264), .Y(
        n20140) );
  nor2_1 U20184 ( .A(n15972), .B(n20111), .Y(n20264) );
  inv_1 U20185 ( .A(n20111), .Y(n20263) );
  o221ai_1 U20186 ( .A1(n20265), .A2(n15920), .B1(n20266), .B2(n18463), .C1(
        n20139), .Y(n20111) );
  nand3_1 U20187 ( .A(n12333), .B(n13401), .C(n12401), .Y(n20139) );
  a21oi_1 U20188 ( .A1(n13307), .A2(n15920), .B1(n20135), .Y(n20266) );
  a21oi_1 U20189 ( .A1(n13307), .A2(n18463), .B1(n20135), .Y(n20265) );
  nand2_1 U20190 ( .A(n20267), .B(n20132), .Y(n20135) );
  nand2_1 U20191 ( .A(n10609), .B(n10775), .Y(n20132) );
  xor2_1 U20192 ( .A(n18532), .B(n20268), .X(n20267) );
  nor2_1 U20193 ( .A(n20129), .B(n20125), .Y(n20268) );
  xnor2_1 U20194 ( .A(n16666), .B(n20269), .Y(n20125) );
  a21oi_1 U20195 ( .A1(n20120), .A2(n12408), .B1(n20270), .Y(n20269) );
  a21oi_1 U20196 ( .A1(n20271), .A2(n15880), .B1(n10608), .Y(n20270) );
  inv_1 U20197 ( .A(n20120), .Y(n20271) );
  xor2_1 U20198 ( .A(n16845), .B(n20272), .X(n20120) );
  a211oi_1 U20199 ( .A1(n12333), .A2(n18455), .B1(n20273), .C1(n20123), .Y(
        n20272) );
  xor2_1 U20200 ( .A(n19960), .B(n20274), .X(n20123) );
  nor2_1 U20201 ( .A(n12331), .B(n24022), .Y(n20274) );
  o21ai_0 U20202 ( .A1(n24022), .A2(n20121), .B1(n17967), .Y(n20273) );
  nor2_1 U20203 ( .A(n24019), .B(n12333), .Y(n20121) );
  xor2_1 U20204 ( .A(n20275), .B(n24045), .X(n20129) );
  nand2_1 U20205 ( .A(n24015), .B(n23993), .Y(n20275) );
  inv_1 U20206 ( .A(n11168), .Y(n18532) );
  o221ai_1 U20207 ( .A1(n24047), .A2(n20276), .B1(n14687), .B2(n14625), .C1(
        n20028), .Y(n11168) );
  inv_1 U20208 ( .A(n20277), .Y(n20028) );
  o21ai_0 U20209 ( .A1(n14702), .A2(n14698), .B1(n19668), .Y(n20277) );
  nand3_1 U20210 ( .A(n14660), .B(n20030), .C(n24047), .Y(n19668) );
  inv_1 U20211 ( .A(n14707), .Y(n14660) );
  nand3_1 U20212 ( .A(n24047), .B(n24046), .C(n24017), .Y(n14625) );
  a222oi_1 U20213 ( .A1(n10636), .A2(n20030), .B1(n14596), .B2(n20252), .C1(
        n14675), .C2(n20033), .Y(n20276) );
  inv_1 U20214 ( .A(n14687), .Y(n14596) );
  nor2_1 U20215 ( .A(n12394), .B(n12305), .Y(n20145) );
  nand4_1 U20216 ( .A(n20278), .B(n20279), .C(n20280), .D(n16182), .Y(n11413)
         );
  nand2_1 U20217 ( .A(n16088), .B(n20281), .Y(n20279) );
  mux2i_1 U20218 ( .A0(n20282), .A1(n20283), .S(n23962), .Y(n20278) );
  nor2_1 U20219 ( .A(n23961), .B(n16170), .Y(n20283) );
  o22ai_1 U20220 ( .A1(n23964), .A2(n16140), .B1(n16087), .B2(n16189), .Y(
        n20282) );
  xnor2_1 U20221 ( .A(n20284), .B(n13307), .Y(n20146) );
  inv_1 U20222 ( .A(n13401), .Y(n13307) );
  nand2_1 U20223 ( .A(n12394), .B(n12305), .Y(n20284) );
  a21oi_1 U20224 ( .A1(n18040), .A2(n20082), .B1(n20080), .Y(n20231) );
  nor2_1 U20225 ( .A(n20082), .B(n18040), .Y(n20080) );
  nand2_1 U20226 ( .A(n12392), .B(n18262), .Y(n20082) );
  inv_1 U20227 ( .A(n16464), .Y(n18040) );
  o221ai_1 U20228 ( .A1(n20285), .A2(n13944), .B1(n24008), .B2(n13951), .C1(
        n13955), .Y(n16464) );
  nand2_1 U20229 ( .A(n13931), .B(n20285), .Y(n13955) );
  xor2_1 U20230 ( .A(n11621), .B(n20286), .X(n20155) );
  nor2_1 U20231 ( .A(n16510), .B(n16545), .Y(n20286) );
  xor2_1 U20232 ( .A(n20287), .B(n18068), .X(n20038) );
  nand2_1 U20233 ( .A(n16545), .B(n16611), .Y(n20287) );
  mux2i_1 U20234 ( .A0(n23986), .A1(n14705), .S(n24042), .Y(n12629) );
  nand3_1 U20235 ( .A(n23922), .B(n10961), .C(n20288), .Y(n10141) );
  mux2i_1 U20236 ( .A0(n20289), .A1(n20290), .S(n23934), .Y(n20288) );
  xor2_1 U20237 ( .A(n10963), .B(n12380), .X(n20290) );
  nor2_1 U20238 ( .A(n10965), .B(n10826), .Y(n20289) );
  nand3_1 U20239 ( .A(n10826), .B(n10964), .C(n10965), .Y(n10961) );
  inv_1 U20240 ( .A(n10963), .Y(n10965) );
  o21ai_0 U20241 ( .A1(n12380), .A2(n20291), .B1(n20292), .Y(n10963) );
  o21ai_0 U20242 ( .A1(n10826), .A2(n20293), .B1(n23935), .Y(n20292) );
  inv_1 U20243 ( .A(n20293), .Y(n20291) );
  inv_1 U20244 ( .A(n23934), .Y(n10964) );
  o22ai_1 U20245 ( .A1(n19449), .A2(n11480), .B1(n11482), .B2(n20294), .Y(
        n10140) );
  xor2_1 U20246 ( .A(n20293), .B(n20295), .X(n20294) );
  xor2_1 U20247 ( .A(n23935), .B(n10826), .X(n20295) );
  o22ai_1 U20248 ( .A1(n16739), .A2(n18747), .B1(n23997), .B2(n20296), .Y(
        n20293) );
  and2_0 U20249 ( .A(n18747), .B(n16739), .X(n20296) );
  o22ai_1 U20250 ( .A1(n11484), .A2(n20297), .B1(n20298), .B2(n20299), .Y(
        n18747) );
  inv_1 U20251 ( .A(n23936), .Y(n20299) );
  nor2_1 U20252 ( .A(n11485), .B(n16744), .Y(n20298) );
  inv_1 U20253 ( .A(n11484), .Y(n16744) );
  inv_1 U20254 ( .A(n11485), .Y(n20297) );
  xor2_1 U20255 ( .A(n20300), .B(n17506), .X(n11485) );
  inv_1 U20256 ( .A(n19466), .Y(n17506) );
  o211ai_1 U20257 ( .A1(n13924), .A2(n19234), .B1(n13946), .C1(n16147), .Y(
        n19466) );
  inv_1 U20258 ( .A(n19239), .Y(n13946) );
  nor2_1 U20259 ( .A(n19745), .B(n13928), .Y(n19239) );
  nand2_1 U20260 ( .A(n23991), .B(n13924), .Y(n19745) );
  o22ai_1 U20261 ( .A1(n16247), .A2(n16248), .B1(n20301), .B2(n16245), .Y(
        n20300) );
  inv_1 U20262 ( .A(n23937), .Y(n16245) );
  and2_0 U20263 ( .A(n16247), .B(n16248), .X(n20301) );
  o21ai_0 U20264 ( .A1(n23950), .A2(n20302), .B1(n20303), .Y(n16248) );
  mux2i_1 U20265 ( .A0(n20304), .A1(n20305), .S(n20306), .Y(n20303) );
  nor2_1 U20266 ( .A(n10607), .B(n20307), .Y(n20305) );
  xor2_1 U20267 ( .A(n20308), .B(n18157), .X(n20302) );
  o22ai_1 U20268 ( .A1(n11665), .A2(n11666), .B1(n20309), .B2(n11667), .Y(
        n16247) );
  inv_1 U20269 ( .A(n70), .Y(n11667) );
  nor2_1 U20270 ( .A(n16325), .B(n20310), .Y(n20309) );
  inv_1 U20271 ( .A(n16325), .Y(n11666) );
  xor2_1 U20272 ( .A(n20311), .B(n20312), .X(n16325) );
  xor2_1 U20273 ( .A(n18163), .B(n20313), .X(n20312) );
  xor2_1 U20274 ( .A(n17860), .B(n23938), .X(n20311) );
  inv_1 U20275 ( .A(n20310), .Y(n11665) );
  o21ai_0 U20276 ( .A1(n23921), .A2(n12929), .B1(n20314), .Y(n20310) );
  xor2_1 U20277 ( .A(n17860), .B(n20315), .X(n20314) );
  nand2_1 U20278 ( .A(n12928), .B(n12930), .Y(n20315) );
  nand2_1 U20279 ( .A(n23921), .B(n12929), .Y(n12930) );
  inv_1 U20280 ( .A(n20316), .Y(n12928) );
  o22ai_1 U20281 ( .A1(n20317), .A2(n16961), .B1(n69), .B2(n20318), .Y(n20316)
         );
  and2_0 U20282 ( .A(n16961), .B(n20317), .X(n20318) );
  o22ai_1 U20283 ( .A1(n16758), .A2(n11404), .B1(n756), .B2(n20319), .Y(n16961) );
  and2_0 U20284 ( .A(n11404), .B(n16758), .X(n20319) );
  xor2_1 U20285 ( .A(n20320), .B(n19327), .X(n11404) );
  o21ai_0 U20286 ( .A1(n12371), .A2(n16295), .B1(n20321), .Y(n20320) );
  xor2_1 U20287 ( .A(n10893), .B(n20322), .X(n20321) );
  o21ai_0 U20288 ( .A1(n11394), .A2(n20323), .B1(n16969), .Y(n20322) );
  o22ai_1 U20289 ( .A1(n16955), .A2(n16608), .B1(n20324), .B2(n10633), .Y(
        n16969) );
  nor2_1 U20290 ( .A(n16762), .B(n20325), .Y(n20324) );
  inv_1 U20291 ( .A(n16955), .Y(n20325) );
  inv_1 U20292 ( .A(n16762), .Y(n16608) );
  xor2_1 U20293 ( .A(n18193), .B(n20326), .X(n16762) );
  xor2_1 U20294 ( .A(n18305), .B(n20327), .X(n20326) );
  xor2_1 U20295 ( .A(n18125), .B(n20328), .X(n16955) );
  a21oi_1 U20296 ( .A1(n11458), .A2(n11460), .B1(n20329), .Y(n20328) );
  inv_1 U20297 ( .A(n20330), .Y(n20329) );
  o21ai_0 U20298 ( .A1(n11460), .A2(n11458), .B1(n23704), .Y(n20330) );
  o22ai_1 U20299 ( .A1(n16233), .A2(n20331), .B1(n23941), .B2(n20332), .Y(
        n11460) );
  nor2_1 U20300 ( .A(n16234), .B(n20333), .Y(n20332) );
  inv_1 U20301 ( .A(n20331), .Y(n16234) );
  o22ai_1 U20302 ( .A1(n16241), .A2(n16240), .B1(n20334), .B2(n11237), .Y(
        n20331) );
  inv_1 U20303 ( .A(n23942), .Y(n11237) );
  and2_0 U20304 ( .A(n16240), .B(n16241), .X(n20334) );
  xnor2_1 U20305 ( .A(n20335), .B(n17385), .Y(n16240) );
  inv_1 U20306 ( .A(n16845), .Y(n17385) );
  o211ai_1 U20307 ( .A1(n11801), .A2(n12357), .B1(n12425), .C1(n20336), .Y(
        n16845) );
  inv_1 U20308 ( .A(n12390), .Y(n12357) );
  nor2_1 U20309 ( .A(n19528), .B(n24033), .Y(n12390) );
  nand2_1 U20310 ( .A(n20337), .B(n11271), .Y(n20335) );
  nand2_1 U20311 ( .A(n23943), .B(n16774), .Y(n11271) );
  xor2_1 U20312 ( .A(n17976), .B(n20338), .X(n20337) );
  nand2_1 U20313 ( .A(n11270), .B(n11268), .Y(n20338) );
  o22ai_1 U20314 ( .A1(n16217), .A2(n16781), .B1(n5), .B2(n20339), .Y(n11268)
         );
  nor2_1 U20315 ( .A(n16216), .B(n20340), .Y(n20339) );
  inv_1 U20316 ( .A(n16781), .Y(n16216) );
  xor2_1 U20317 ( .A(n20341), .B(n20342), .X(n16781) );
  xor2_1 U20318 ( .A(n18320), .B(n20343), .X(n20342) );
  xor2_1 U20319 ( .A(n15902), .B(n12297), .X(n20341) );
  inv_1 U20320 ( .A(n20340), .Y(n16217) );
  o21ai_0 U20321 ( .A1(n11218), .A2(n7), .B1(n11217), .Y(n20340) );
  nand2_1 U20322 ( .A(n16785), .B(n20344), .Y(n11217) );
  nor2_1 U20323 ( .A(n20344), .B(n16785), .Y(n11218) );
  xnor2_1 U20324 ( .A(n18390), .B(n20345), .Y(n16785) );
  xor2_1 U20325 ( .A(n10606), .B(n20346), .X(n20345) );
  o22ai_1 U20326 ( .A1(n11295), .A2(n16788), .B1(n23945), .B2(n20347), .Y(
        n20344) );
  nor2_1 U20327 ( .A(n11296), .B(n20348), .Y(n20347) );
  inv_1 U20328 ( .A(n11295), .Y(n20348) );
  inv_1 U20329 ( .A(n16788), .Y(n11296) );
  xor2_1 U20330 ( .A(n20349), .B(n20350), .X(n16788) );
  xor2_1 U20331 ( .A(n20351), .B(n11209), .X(n11295) );
  inv_1 U20332 ( .A(n18125), .Y(n11209) );
  o22ai_1 U20333 ( .A1(n16211), .A2(n20352), .B1(n23909), .B2(n20353), .Y(
        n20351) );
  nor2_1 U20334 ( .A(n16209), .B(n16791), .Y(n20353) );
  inv_1 U20335 ( .A(n16209), .Y(n20352) );
  xnor2_1 U20336 ( .A(n20354), .B(n17774), .Y(n16209) );
  nand3_1 U20337 ( .A(n20355), .B(n20088), .C(n20356), .Y(n17774) );
  a221oi_1 U20338 ( .A1(n23976), .A2(n20357), .B1(n16107), .B2(n20093), .C1(
        n19408), .Y(n20356) );
  inv_1 U20339 ( .A(n19951), .Y(n19408) );
  inv_1 U20340 ( .A(n16164), .Y(n20093) );
  o21ai_0 U20341 ( .A1(n23975), .A2(n23977), .B1(n20358), .Y(n20357) );
  inv_1 U20342 ( .A(n20359), .Y(n20088) );
  o22ai_1 U20343 ( .A1(n16124), .A2(n16178), .B1(n19407), .B2(n16154), .Y(
        n20359) );
  nand2_1 U20344 ( .A(n19955), .B(n16163), .Y(n16154) );
  mux2i_1 U20345 ( .A0(n16173), .A1(n20360), .S(n23978), .Y(n20355) );
  o22ai_1 U20346 ( .A1(n20361), .A2(n12519), .B1(n20362), .B2(n11197), .Y(
        n20354) );
  inv_1 U20347 ( .A(n23946), .Y(n11197) );
  nor2_1 U20348 ( .A(n12523), .B(n16495), .Y(n20362) );
  inv_1 U20349 ( .A(n12519), .Y(n16495) );
  inv_1 U20350 ( .A(n20361), .Y(n12523) );
  o21ai_0 U20351 ( .A1(n23981), .A2(n20363), .B1(n20364), .Y(n12519) );
  mux2i_1 U20352 ( .A0(n20365), .A1(n20366), .S(n20367), .Y(n20364) );
  nor2_1 U20353 ( .A(n18303), .B(n15999), .Y(n20366) );
  xor2_1 U20354 ( .A(n20368), .B(n18400), .X(n20363) );
  o21ai_0 U20355 ( .A1(n16643), .A2(n12735), .B1(n20369), .Y(n20361) );
  xor2_1 U20356 ( .A(n17232), .B(n20370), .X(n20369) );
  nor2_1 U20357 ( .A(n11156), .B(n11153), .Y(n20370) );
  o221ai_1 U20358 ( .A1(n698), .A2(n20371), .B1(n12469), .B2(n20372), .C1(
        n20373), .Y(n11153) );
  nand2_1 U20359 ( .A(n12470), .B(n11489), .Y(n20373) );
  xor2_1 U20360 ( .A(n12632), .B(n10638), .X(n12470) );
  inv_1 U20361 ( .A(n12632), .Y(n20372) );
  inv_1 U20362 ( .A(n20374), .Y(n12469) );
  a21oi_1 U20363 ( .A1(n12632), .A2(n11751), .B1(n20374), .Y(n20371) );
  o22ai_1 U20364 ( .A1(n20375), .A2(n12745), .B1(n52), .B2(n20376), .Y(n20374)
         );
  nor2_1 U20365 ( .A(n20377), .B(n12744), .Y(n20376) );
  inv_1 U20366 ( .A(n20375), .Y(n12744) );
  inv_1 U20367 ( .A(n12745), .Y(n20377) );
  xor2_1 U20368 ( .A(n20378), .B(n18066), .X(n12745) );
  nor2_1 U20369 ( .A(n20379), .B(n13833), .Y(n18066) );
  nor3_1 U20370 ( .A(n10624), .B(n24008), .C(n13951), .Y(n13833) );
  mux2i_1 U20371 ( .A0(n13956), .A1(n13943), .S(n24009), .Y(n20379) );
  o22ai_1 U20372 ( .A1(n11347), .A2(n11348), .B1(n54), .B2(n20380), .Y(n20378)
         );
  and2_0 U20373 ( .A(n11348), .B(n11347), .X(n20380) );
  xnor2_1 U20374 ( .A(n20381), .B(n11103), .Y(n11348) );
  a211oi_1 U20375 ( .A1(n13944), .A2(n20285), .B1(n20382), .C1(n13860), .Y(
        n11103) );
  nor2_1 U20376 ( .A(n18668), .B(n13944), .Y(n13860) );
  o22ai_1 U20377 ( .A1(n11550), .A2(n11548), .B1(n20383), .B2(n20384), .Y(
        n20381) );
  inv_1 U20378 ( .A(n23969), .Y(n20384) );
  and2_0 U20379 ( .A(n11548), .B(n11550), .X(n20383) );
  xor2_1 U20380 ( .A(n20385), .B(n20386), .X(n11548) );
  nand2_1 U20381 ( .A(n20387), .B(n20388), .Y(n20385) );
  a21oi_1 U20382 ( .A1(n17021), .A2(n16799), .B1(n20389), .Y(n11550) );
  xor2_1 U20383 ( .A(n10919), .B(n20390), .X(n20389) );
  nor2_1 U20384 ( .A(n17022), .B(n17020), .Y(n20390) );
  o22ai_1 U20385 ( .A1(n16804), .A2(n17027), .B1(n23925), .B2(n20391), .Y(
        n17020) );
  and2_0 U20386 ( .A(n17027), .B(n16804), .X(n20391) );
  o21ai_0 U20387 ( .A1(n23706), .A2(n16198), .B1(n20392), .Y(n17027) );
  xor2_1 U20388 ( .A(n12806), .B(n20393), .X(n20392) );
  a21oi_1 U20389 ( .A1(n23706), .A2(n16198), .B1(n11568), .Y(n20393) );
  o22ai_1 U20390 ( .A1(n11778), .A2(n20394), .B1(n20395), .B2(n20396), .Y(
        n11568) );
  inv_1 U20391 ( .A(n23971), .Y(n20396) );
  nor2_1 U20392 ( .A(n10777), .B(n12807), .Y(n20395) );
  inv_1 U20393 ( .A(n10777), .Y(n20394) );
  xor2_1 U20394 ( .A(n20397), .B(n20398), .X(n10777) );
  xor2_1 U20395 ( .A(n15913), .B(n16246), .X(n20398) );
  inv_1 U20396 ( .A(n17737), .Y(n16246) );
  a221oi_1 U20397 ( .A1(n13944), .A2(n20382), .B1(n24009), .B2(n13845), .C1(
        n13862), .Y(n17737) );
  inv_1 U20398 ( .A(n13764), .Y(n13862) );
  nor2_1 U20399 ( .A(n13943), .B(n13940), .Y(n20382) );
  inv_1 U20400 ( .A(n13939), .Y(n13943) );
  xor2_1 U20401 ( .A(n18432), .B(n20399), .X(n20397) );
  inv_1 U20402 ( .A(n12807), .Y(n11778) );
  nand2_1 U20403 ( .A(n12521), .B(n11779), .Y(n12807) );
  xor2_1 U20404 ( .A(n18284), .B(n20400), .X(n11779) );
  xor2_1 U20405 ( .A(n15920), .B(n20401), .X(n20400) );
  a21oi_1 U20406 ( .A1(n24013), .A2(n18672), .B1(n13341), .Y(n12806) );
  nor2_1 U20407 ( .A(n13399), .B(n23983), .Y(n13341) );
  inv_1 U20408 ( .A(n13379), .Y(n18672) );
  inv_1 U20409 ( .A(n16197), .Y(n16198) );
  xor2_1 U20410 ( .A(n20402), .B(n20403), .X(n16197) );
  xor2_1 U20411 ( .A(n20404), .B(n24011), .X(n20402) );
  xnor2_1 U20412 ( .A(n20405), .B(n20406), .Y(n16804) );
  xor2_1 U20413 ( .A(n20407), .B(n18292), .X(n20406) );
  xor2_1 U20414 ( .A(n20408), .B(n19507), .X(n20405) );
  inv_1 U20415 ( .A(n18840), .Y(n19507) );
  xor2_1 U20416 ( .A(n11622), .B(n23993), .X(n20408) );
  o211ai_1 U20417 ( .A1(n13957), .A2(n19234), .B1(n16147), .C1(n13962), .Y(
        n11622) );
  inv_1 U20418 ( .A(n19856), .Y(n13962) );
  nor2_1 U20419 ( .A(n13930), .B(n19235), .Y(n19856) );
  nor2_1 U20420 ( .A(n17021), .B(n16799), .Y(n17022) );
  xor2_1 U20421 ( .A(n20409), .B(n18420), .X(n16799) );
  xor2_1 U20422 ( .A(n20410), .B(n12401), .X(n20409) );
  inv_1 U20423 ( .A(n23924), .Y(n17021) );
  xor2_1 U20424 ( .A(n20411), .B(n20412), .X(n11347) );
  xor2_1 U20425 ( .A(n12388), .B(n11710), .X(n20412) );
  xor2_1 U20426 ( .A(n20413), .B(n18409), .X(n20411) );
  xor2_1 U20427 ( .A(n20414), .B(n18417), .X(n20375) );
  inv_1 U20428 ( .A(n18411), .Y(n18417) );
  nand2_1 U20429 ( .A(n20415), .B(n20416), .Y(n20414) );
  inv_1 U20430 ( .A(n11489), .Y(n11751) );
  xor2_1 U20431 ( .A(n20417), .B(n20418), .X(n12632) );
  xor2_1 U20432 ( .A(n23987), .B(n20419), .X(n20418) );
  xor2_1 U20433 ( .A(n20420), .B(n18999), .X(n20417) );
  nor2_1 U20434 ( .A(n11155), .B(n12473), .Y(n11156) );
  inv_1 U20435 ( .A(n16643), .Y(n11155) );
  inv_1 U20436 ( .A(n11159), .Y(n17232) );
  o221ai_1 U20437 ( .A1(n23992), .A2(n13930), .B1(n19235), .B2(n19236), .C1(
        n20421), .Y(n11159) );
  mux2i_1 U20438 ( .A0(n19747), .A1(n13924), .S(n13938), .Y(n20421) );
  inv_1 U20439 ( .A(n12473), .Y(n12735) );
  xor2_1 U20440 ( .A(n20422), .B(n20423), .X(n16643) );
  xor2_1 U20441 ( .A(n18223), .B(n12394), .X(n20422) );
  inv_1 U20442 ( .A(n16791), .Y(n16211) );
  o21ai_0 U20443 ( .A1(n15990), .A2(n20424), .B1(n20425), .Y(n16791) );
  mux2i_1 U20444 ( .A0(n20426), .A1(n20427), .S(n20428), .Y(n20425) );
  nor2_1 U20445 ( .A(n12392), .B(n18309), .Y(n20427) );
  xor2_1 U20446 ( .A(n20428), .B(n18309), .X(n20424) );
  or2_0 U20447 ( .A(n16774), .B(n23943), .X(n11270) );
  xor2_1 U20448 ( .A(n20429), .B(n18382), .X(n16774) );
  xor2_1 U20449 ( .A(n20430), .B(n23958), .X(n20429) );
  xor2_1 U20450 ( .A(n20431), .B(n20432), .X(n16241) );
  xor2_1 U20451 ( .A(n19960), .B(n20433), .X(n20432) );
  xor2_1 U20452 ( .A(n16545), .B(n24045), .X(n20433) );
  nand2_1 U20453 ( .A(n20434), .B(n13377), .Y(n19960) );
  nand3_1 U20454 ( .A(n24003), .B(n19562), .C(n24020), .Y(n13377) );
  mux2i_1 U20455 ( .A0(n13387), .A1(n13385), .S(n24020), .Y(n20434) );
  xor2_1 U20456 ( .A(n18371), .B(n20435), .X(n20431) );
  inv_1 U20457 ( .A(n20333), .Y(n16233) );
  o21ai_0 U20458 ( .A1(n20436), .A2(n16524), .B1(n20437), .Y(n20333) );
  mux2i_1 U20459 ( .A0(n20438), .A1(n20439), .S(n20440), .Y(n20437) );
  nor2_1 U20460 ( .A(n12319), .B(n18377), .Y(n20439) );
  xor2_1 U20461 ( .A(n20441), .B(n18373), .X(n20436) );
  o21ai_0 U20462 ( .A1(n20442), .A2(n15931), .B1(n20443), .Y(n11458) );
  mux2i_1 U20463 ( .A0(n20444), .A1(n20445), .S(n20446), .Y(n20443) );
  nor2_1 U20464 ( .A(n12302), .B(n18336), .Y(n20445) );
  xor2_1 U20465 ( .A(n18336), .B(n20446), .X(n20442) );
  o221ai_1 U20466 ( .A1(n24025), .A2(n12385), .B1(n12223), .B2(n12334), .C1(
        n20187), .Y(n18125) );
  a21oi_1 U20467 ( .A1(n20258), .A2(n20447), .B1(n19684), .Y(n20187) );
  inv_1 U20468 ( .A(n16295), .Y(n20323) );
  inv_1 U20469 ( .A(n12371), .Y(n11394) );
  o221ai_1 U20470 ( .A1(n13928), .A2(n13950), .B1(n23991), .B2(n13957), .C1(
        n19234), .Y(n10893) );
  xor2_1 U20471 ( .A(n20448), .B(n18192), .X(n16295) );
  xor2_1 U20472 ( .A(n16611), .B(n20449), .X(n20448) );
  inv_1 U20473 ( .A(n11405), .Y(n16758) );
  o21ai_0 U20474 ( .A1(n12299), .A2(n20450), .B1(n20451), .Y(n11405) );
  mux2i_1 U20475 ( .A0(n20452), .A1(n20453), .S(n20454), .Y(n20451) );
  nor2_1 U20476 ( .A(n18346), .B(n15955), .Y(n20453) );
  xor2_1 U20477 ( .A(n20455), .B(n18181), .X(n20450) );
  inv_1 U20478 ( .A(n16752), .Y(n20317) );
  xor2_1 U20479 ( .A(n20456), .B(n20457), .X(n16752) );
  xor2_1 U20480 ( .A(n20458), .B(n18178), .X(n20457) );
  xor2_1 U20481 ( .A(n17746), .B(n23951), .X(n20456) );
  o211ai_1 U20482 ( .A1(n18845), .A2(n16176), .B1(n20459), .C1(n20460), .Y(
        n17746) );
  a221oi_1 U20483 ( .A1(n23976), .A2(n16134), .B1(n16173), .B2(n16071), .C1(
        n18844), .Y(n20460) );
  nor2_1 U20484 ( .A(n16121), .B(n19407), .Y(n18844) );
  nand2_1 U20485 ( .A(n23975), .B(n19415), .Y(n16121) );
  mux2i_1 U20486 ( .A0(n20461), .A1(n20462), .S(n23977), .Y(n20459) );
  o21ai_0 U20487 ( .A1(n16163), .A2(n16164), .B1(n16188), .Y(n20461) );
  o21ai_0 U20488 ( .A1(n24020), .A2(n19560), .B1(n13164), .Y(n17860) );
  nand3_1 U20489 ( .A(n24003), .B(n13385), .C(n24020), .Y(n13164) );
  xor2_1 U20490 ( .A(n20463), .B(n20464), .X(n12929) );
  xor2_1 U20491 ( .A(n15953), .B(n17152), .X(n20464) );
  nand4_1 U20492 ( .A(n20465), .B(n12404), .C(n12396), .D(n12385), .Y(n17152)
         );
  nand2_1 U20493 ( .A(n24025), .B(n24035), .Y(n12396) );
  nand2_1 U20494 ( .A(n12422), .B(n24025), .Y(n20465) );
  xor2_1 U20495 ( .A(n20466), .B(n18166), .X(n20463) );
  xor2_1 U20496 ( .A(n20188), .B(n20467), .X(n11484) );
  a21oi_1 U20497 ( .A1(n18764), .A2(n20467), .B1(n18765), .Y(n16739) );
  inv_1 U20498 ( .A(n20468), .Y(n20467) );
  o22ai_1 U20499 ( .A1(n23950), .A2(n20307), .B1(n20306), .B2(n20469), .Y(
        n20468) );
  xor2_1 U20500 ( .A(n18947), .B(n20304), .X(n20469) );
  nor2_1 U20501 ( .A(n10607), .B(n18157), .Y(n20304) );
  nand4_1 U20502 ( .A(n20470), .B(n13907), .C(n13764), .D(n16146), .Y(n18947)
         );
  nand2_1 U20503 ( .A(n1678), .B(n18443), .Y(n16146) );
  nor2_1 U20504 ( .A(n13944), .B(n24008), .Y(n18443) );
  nand2_1 U20505 ( .A(n13940), .B(n20285), .Y(n13764) );
  inv_1 U20506 ( .A(n13956), .Y(n20285) );
  nand2_1 U20507 ( .A(n24008), .B(n10624), .Y(n13956) );
  nand2_1 U20508 ( .A(n13844), .B(n13939), .Y(n13907) );
  inv_1 U20509 ( .A(n18445), .Y(n13844) );
  nand2_1 U20510 ( .A(n23972), .B(n10626), .Y(n18445) );
  nand3_1 U20511 ( .A(n13951), .B(n13944), .C(n13845), .Y(n20470) );
  inv_1 U20512 ( .A(n18668), .Y(n13845) );
  nand2_1 U20513 ( .A(n24009), .B(n23972), .Y(n13944) );
  inv_1 U20514 ( .A(n20308), .Y(n20306) );
  o221ai_1 U20515 ( .A1(n20471), .A2(n16013), .B1(n18163), .B2(n20313), .C1(
        n20472), .Y(n20308) );
  o21ai_0 U20516 ( .A1(n18163), .A2(n16013), .B1(n17550), .Y(n20472) );
  inv_1 U20517 ( .A(n20473), .Y(n20471) );
  o21ai_0 U20518 ( .A1(n17550), .A2(n18163), .B1(n20313), .Y(n20473) );
  xor2_1 U20519 ( .A(n20474), .B(n18999), .X(n20313) );
  o22ai_1 U20520 ( .A1(n18350), .A2(n20475), .B1(n20476), .B2(n15953), .Y(
        n20474) );
  nor2_1 U20521 ( .A(n20466), .B(n18166), .Y(n20476) );
  inv_1 U20522 ( .A(n18350), .Y(n18166) );
  inv_1 U20523 ( .A(n20466), .Y(n20475) );
  xor2_1 U20524 ( .A(n20477), .B(n19382), .X(n20466) );
  inv_1 U20525 ( .A(n17573), .Y(n19382) );
  nand4_1 U20526 ( .A(n20478), .B(n20479), .C(n20280), .D(n16186), .Y(n17573)
         );
  nand2_1 U20527 ( .A(n16162), .B(n16088), .Y(n16186) );
  inv_1 U20528 ( .A(n16144), .Y(n16088) );
  nand3_1 U20529 ( .A(n23962), .B(n10616), .C(n16162), .Y(n20280) );
  inv_1 U20530 ( .A(n16180), .Y(n16162) );
  nand2_1 U20531 ( .A(n20480), .B(n20281), .Y(n16180) );
  nand2_1 U20532 ( .A(n16137), .B(n16168), .Y(n20479) );
  inv_1 U20533 ( .A(n16170), .Y(n16168) );
  nand2_1 U20534 ( .A(n23960), .B(n23963), .Y(n16170) );
  mux2i_1 U20535 ( .A0(n20481), .A1(n20482), .S(n23962), .Y(n20478) );
  mux2i_1 U20536 ( .A0(n16144), .A1(n16179), .S(n23963), .Y(n20482) );
  nand2_1 U20537 ( .A(n10616), .B(n20046), .Y(n16144) );
  inv_1 U20538 ( .A(n23961), .Y(n20046) );
  nand3_1 U20539 ( .A(n16191), .B(n14215), .C(n16182), .Y(n20481) );
  nand2_1 U20540 ( .A(n16172), .B(n16100), .Y(n16182) );
  inv_1 U20541 ( .A(n16189), .Y(n16172) );
  nand2_1 U20542 ( .A(n16087), .B(n20051), .Y(n14215) );
  inv_1 U20543 ( .A(n16179), .Y(n20051) );
  nand2_1 U20544 ( .A(n23961), .B(n10616), .Y(n16179) );
  nand2_1 U20545 ( .A(n16101), .B(n16087), .Y(n16191) );
  o22ai_1 U20546 ( .A1(n18178), .A2(n20458), .B1(n20483), .B2(n20209), .Y(
        n20477) );
  and2_0 U20547 ( .A(n20458), .B(n18178), .X(n20483) );
  o21ai_0 U20548 ( .A1(n12299), .A2(n18346), .B1(n20484), .Y(n20458) );
  xor2_1 U20549 ( .A(n20485), .B(n10928), .X(n20484) );
  inv_1 U20550 ( .A(n11677), .Y(n10928) );
  o22ai_1 U20551 ( .A1(n20068), .A2(n13381), .B1(n20486), .B2(n13403), .Y(
        n11677) );
  or2_0 U20552 ( .A(n20454), .B(n20452), .X(n20485) );
  nor2_1 U20553 ( .A(n18181), .B(n15955), .Y(n20452) );
  inv_1 U20554 ( .A(n18346), .Y(n18181) );
  inv_1 U20555 ( .A(n20455), .Y(n20454) );
  o22ai_1 U20556 ( .A1(n18345), .A2(n20487), .B1(n20488), .B2(n16611), .Y(
        n20455) );
  nor2_1 U20557 ( .A(n20449), .B(n18192), .Y(n20488) );
  inv_1 U20558 ( .A(n18345), .Y(n18192) );
  inv_1 U20559 ( .A(n20487), .Y(n20449) );
  o22ai_1 U20560 ( .A1(n18193), .A2(n20327), .B1(n20489), .B2(n18305), .Y(
        n20487) );
  inv_1 U20561 ( .A(n23948), .Y(n18305) );
  and2_0 U20562 ( .A(n20327), .B(n18193), .X(n20489) );
  nand2_1 U20563 ( .A(n20490), .B(n20491), .Y(n20327) );
  xor2_1 U20564 ( .A(n10946), .B(n20492), .X(n20491) );
  nor2_1 U20565 ( .A(n18336), .B(n15931), .Y(n20492) );
  inv_1 U20566 ( .A(n16848), .Y(n10946) );
  nand3_1 U20567 ( .A(n20493), .B(n19862), .C(n20494), .Y(n16848) );
  nor3_1 U20568 ( .A(n12329), .B(n11822), .C(n20495), .Y(n20494) );
  inv_1 U20569 ( .A(n20013), .Y(n20495) );
  nand3_1 U20570 ( .A(n12407), .B(n20496), .C(n20007), .Y(n20013) );
  inv_1 U20571 ( .A(n24027), .Y(n12407) );
  nor2_1 U20572 ( .A(n20021), .B(n24029), .Y(n11822) );
  inv_1 U20573 ( .A(n19865), .Y(n20021) );
  nor2_1 U20574 ( .A(n12416), .B(n24024), .Y(n19865) );
  nor2_1 U20575 ( .A(n10610), .B(n20005), .Y(n12329) );
  or2_0 U20576 ( .A(n12370), .B(n24024), .X(n20005) );
  nand2_1 U20577 ( .A(n20016), .B(n20007), .Y(n19862) );
  inv_1 U20578 ( .A(n12428), .Y(n20016) );
  nand2_1 U20579 ( .A(n24030), .B(n12387), .Y(n12428) );
  mux2i_1 U20580 ( .A0(n20497), .A1(n20498), .S(n24027), .Y(n20493) );
  o21ai_0 U20581 ( .A1(n20496), .A2(n12374), .B1(n20245), .Y(n20498) );
  nand2_1 U20582 ( .A(n19864), .B(n20496), .Y(n20245) );
  inv_1 U20583 ( .A(n19315), .Y(n19864) );
  nand3_1 U20584 ( .A(n24028), .B(n10610), .C(n24024), .Y(n19315) );
  o21ai_0 U20585 ( .A1(n20007), .A2(n12416), .B1(n12370), .Y(n20497) );
  nand2_1 U20586 ( .A(n12387), .B(n20496), .Y(n12370) );
  inv_1 U20587 ( .A(n24030), .Y(n20496) );
  inv_1 U20588 ( .A(n24028), .Y(n12387) );
  nand2_1 U20589 ( .A(n24030), .B(n24028), .Y(n12416) );
  inv_1 U20590 ( .A(n12374), .Y(n20007) );
  nand2_1 U20591 ( .A(n24029), .B(n24024), .Y(n12374) );
  xnor2_1 U20592 ( .A(n11292), .B(n20499), .Y(n20490) );
  nor2_1 U20593 ( .A(n20444), .B(n20446), .Y(n20499) );
  a21oi_1 U20594 ( .A1(n18373), .A2(n12319), .B1(n20500), .Y(n20446) );
  xor2_1 U20595 ( .A(n18118), .B(n20501), .X(n20500) );
  or2_0 U20596 ( .A(n20440), .B(n20438), .X(n20501) );
  nor2_1 U20597 ( .A(n18373), .B(n12319), .Y(n20438) );
  inv_1 U20598 ( .A(n20441), .Y(n20440) );
  o221ai_1 U20599 ( .A1(n20502), .A2(n16545), .B1(n18329), .B2(n20503), .C1(
        n20504), .Y(n20441) );
  o21ai_0 U20600 ( .A1(n16545), .A2(n18329), .B1(n17611), .Y(n20504) );
  inv_1 U20601 ( .A(n18371), .Y(n18329) );
  inv_1 U20602 ( .A(n23959), .Y(n16545) );
  a21oi_1 U20603 ( .A1(n18371), .A2(n18397), .B1(n20435), .Y(n20502) );
  inv_1 U20604 ( .A(n20503), .Y(n20435) );
  o22ai_1 U20605 ( .A1(n20505), .A2(n18382), .B1(n20506), .B2(n18413), .Y(
        n20503) );
  nor2_1 U20606 ( .A(n18386), .B(n20430), .Y(n20506) );
  inv_1 U20607 ( .A(n18382), .Y(n18386) );
  xnor2_1 U20608 ( .A(n20507), .B(n20508), .Y(n18382) );
  inv_1 U20609 ( .A(n20430), .Y(n20505) );
  o22ai_1 U20610 ( .A1(n18320), .A2(n20343), .B1(n20509), .B2(n15902), .Y(
        n20430) );
  and2_0 U20611 ( .A(n18320), .B(n20343), .X(n20509) );
  xnor2_1 U20612 ( .A(n14685), .B(n20510), .Y(n20343) );
  a21oi_1 U20613 ( .A1(n20511), .A2(n18315), .B1(n20512), .Y(n20510) );
  a21oi_1 U20614 ( .A1(n18390), .A2(n20346), .B1(n10606), .Y(n20512) );
  inv_1 U20615 ( .A(n18390), .Y(n18315) );
  xor2_1 U20616 ( .A(n20513), .B(n20514), .X(n18390) );
  xor2_1 U20617 ( .A(n23959), .B(n12393), .X(n20514) );
  inv_1 U20618 ( .A(n20346), .Y(n20511) );
  o221ai_1 U20619 ( .A1(n18394), .A2(n20349), .B1(n10920), .B2(n20350), .C1(
        n20515), .Y(n20346) );
  o21ai_0 U20620 ( .A1(n20516), .A2(n20517), .B1(n16510), .Y(n20515) );
  inv_1 U20621 ( .A(n20349), .Y(n20517) );
  nor2_1 U20622 ( .A(n18394), .B(n17066), .Y(n20516) );
  xor2_1 U20623 ( .A(n18311), .B(n12340), .X(n20350) );
  inv_1 U20624 ( .A(n17066), .Y(n10920) );
  o211ai_1 U20625 ( .A1(n12423), .A2(n19529), .B1(n12425), .C1(n20518), .Y(
        n17066) );
  mux2i_1 U20626 ( .A0(n19531), .A1(n19875), .S(n12384), .Y(n20518) );
  inv_1 U20627 ( .A(n12405), .Y(n19875) );
  o21ai_0 U20628 ( .A1(n15990), .A2(n18309), .B1(n20519), .Y(n20349) );
  xor2_1 U20629 ( .A(n16750), .B(n20520), .X(n20519) );
  nor2_1 U20630 ( .A(n20426), .B(n20428), .Y(n20520) );
  a21oi_1 U20631 ( .A1(n15999), .A2(n18400), .B1(n20521), .Y(n20428) );
  xor2_1 U20632 ( .A(n20522), .B(n17958), .X(n20521) );
  inv_1 U20633 ( .A(n16868), .Y(n17958) );
  mux2i_1 U20634 ( .A0(n14697), .A1(n14666), .S(n24042), .Y(n16868) );
  inv_1 U20635 ( .A(n14661), .Y(n14666) );
  nand2_1 U20636 ( .A(n24040), .B(n23986), .Y(n14697) );
  or2_0 U20637 ( .A(n20367), .B(n20365), .X(n20522) );
  nor2_1 U20638 ( .A(n18400), .B(n15999), .Y(n20365) );
  inv_1 U20639 ( .A(n20368), .Y(n20367) );
  o22ai_1 U20640 ( .A1(n18222), .A2(n20423), .B1(n20523), .B2(n15992), .Y(
        n20368) );
  nor2_1 U20641 ( .A(n18223), .B(n20524), .Y(n20523) );
  inv_1 U20642 ( .A(n20524), .Y(n20423) );
  o22ai_1 U20643 ( .A1(n20420), .A2(n16453), .B1(n20419), .B2(n20525), .Y(
        n20524) );
  xor2_1 U20644 ( .A(n12823), .B(n20526), .X(n20525) );
  nor2_1 U20645 ( .A(n23987), .B(n18406), .Y(n20526) );
  inv_1 U20646 ( .A(n20420), .Y(n18406) );
  inv_1 U20647 ( .A(n18052), .Y(n12823) );
  nor2_1 U20648 ( .A(n20527), .B(n20528), .Y(n18052) );
  mux2i_1 U20649 ( .A0(n13403), .A1(n13379), .S(n20529), .Y(n20527) );
  a21oi_1 U20650 ( .A1(n20415), .A2(n18411), .B1(n20530), .Y(n20419) );
  inv_1 U20651 ( .A(n20416), .Y(n20530) );
  o221ai_1 U20652 ( .A1(n12388), .A2(n20531), .B1(n18409), .B2(n20532), .C1(
        n18262), .Y(n20416) );
  nor2_1 U20653 ( .A(n18296), .B(n20413), .Y(n20531) );
  xor2_1 U20654 ( .A(n20533), .B(n20534), .X(n18411) );
  xor2_1 U20655 ( .A(n18405), .B(n16000), .X(n20534) );
  o21ai_0 U20656 ( .A1(n23987), .A2(n15999), .B1(n16001), .Y(n16000) );
  nand2_1 U20657 ( .A(n23987), .B(n15999), .Y(n16001) );
  inv_1 U20658 ( .A(n11301), .Y(n18405) );
  a221oi_1 U20659 ( .A1(n13379), .A2(n20068), .B1(n23983), .B2(n18673), .C1(
        n20535), .Y(n11301) );
  o21ai_0 U20660 ( .A1(n13403), .A2(n24013), .B1(n20536), .Y(n20535) );
  inv_1 U20661 ( .A(n13399), .Y(n18673) );
  nand2_1 U20662 ( .A(n23983), .B(n23982), .Y(n13379) );
  o211ai_1 U20663 ( .A1(n18296), .A2(n20413), .B1(n20537), .C1(n23985), .Y(
        n20415) );
  o21ai_0 U20664 ( .A1(n18409), .A2(n20532), .B1(n12388), .Y(n20537) );
  inv_1 U20665 ( .A(n20413), .Y(n20532) );
  inv_1 U20666 ( .A(n18296), .Y(n18409) );
  xnor2_1 U20667 ( .A(n20538), .B(n12686), .Y(n20413) );
  nand3_1 U20668 ( .A(n13399), .B(n13392), .C(n20539), .Y(n12686) );
  a22oi_1 U20669 ( .A1(n24012), .A2(n13398), .B1(n20068), .B2(n10622), .Y(
        n20539) );
  nand2_1 U20670 ( .A(n20486), .B(n23982), .Y(n13399) );
  inv_1 U20671 ( .A(n13404), .Y(n20486) );
  nand2_1 U20672 ( .A(n24012), .B(n18468), .Y(n13404) );
  nand2_1 U20673 ( .A(n20540), .B(n20388), .Y(n20538) );
  nand2_1 U20674 ( .A(n18293), .B(n12305), .Y(n20388) );
  xor2_1 U20675 ( .A(n11574), .B(n20541), .X(n20540) );
  nand2_1 U20676 ( .A(n20386), .B(n20542), .Y(n20541) );
  xnor2_1 U20677 ( .A(n20387), .B(n11048), .Y(n20542) );
  mux2i_1 U20678 ( .A0(n20543), .A1(n16181), .S(n10605), .Y(n11048) );
  or2_0 U20679 ( .A(n18293), .B(n12305), .X(n20387) );
  xnor2_1 U20680 ( .A(n20544), .B(n20545), .Y(n18293) );
  xor2_1 U20681 ( .A(n16931), .B(n20546), .X(n20545) );
  inv_1 U20682 ( .A(n20547), .Y(n20386) );
  o22ai_1 U20683 ( .A1(n18241), .A2(n20410), .B1(n20548), .B2(n18463), .Y(
        n20547) );
  and2_0 U20684 ( .A(n20410), .B(n18241), .X(n20548) );
  o22ai_1 U20685 ( .A1(n18292), .A2(n20407), .B1(n20549), .B2(n10775), .Y(
        n20410) );
  and2_0 U20686 ( .A(n20407), .B(n18292), .X(n20549) );
  o22ai_1 U20687 ( .A1(n20403), .A2(n20404), .B1(n24011), .B2(n20550), .Y(
        n20407) );
  and2_0 U20688 ( .A(n20404), .B(n20403), .X(n20550) );
  o22ai_1 U20689 ( .A1(n18432), .A2(n15913), .B1(n20399), .B2(n20551), .Y(
        n20404) );
  xor2_1 U20690 ( .A(n18379), .B(n20552), .X(n20551) );
  nor2_1 U20691 ( .A(n24022), .B(n18429), .Y(n20552) );
  inv_1 U20692 ( .A(n18432), .Y(n18429) );
  nand4_1 U20693 ( .A(n19951), .B(n16178), .C(n20553), .D(n20554), .Y(n18379)
         );
  a222oi_1 U20694 ( .A1(n16124), .A2(n19415), .B1(n16173), .B2(n16071), .C1(
        n23974), .C2(n16134), .Y(n20554) );
  nor2_1 U20695 ( .A(n16164), .B(n23975), .Y(n16173) );
  a22oi_1 U20696 ( .A1(n16113), .A2(n23978), .B1(n16107), .B2(n16053), .Y(
        n20553) );
  inv_1 U20697 ( .A(n16139), .Y(n16053) );
  nand2_1 U20698 ( .A(n19411), .B(n19415), .Y(n16139) );
  nor2_1 U20699 ( .A(n23974), .B(n23975), .Y(n19411) );
  nor2_1 U20700 ( .A(n23978), .B(n23977), .Y(n16107) );
  nand2_1 U20701 ( .A(n16113), .B(n23977), .Y(n19951) );
  nor2_1 U20702 ( .A(n20092), .B(n16163), .Y(n16113) );
  a22oi_1 U20703 ( .A1(n20401), .A2(n18284), .B1(n15920), .B2(n20555), .Y(
        n20399) );
  or2_0 U20704 ( .A(n18284), .B(n20401), .X(n20555) );
  xor2_1 U20705 ( .A(n20556), .B(n20557), .X(n18284) );
  xor2_1 U20706 ( .A(n20558), .B(n18136), .X(n20556) );
  a221oi_1 U20707 ( .A1(n10626), .A2(n13939), .B1(n24008), .B2(n13931), .C1(
        n18444), .Y(n18136) );
  o22ai_1 U20708 ( .A1(n24008), .A2(n13951), .B1(n10626), .B2(n18668), .Y(
        n18444) );
  nand2_1 U20709 ( .A(n24008), .B(n1678), .Y(n18668) );
  inv_1 U20710 ( .A(n13940), .Y(n13951) );
  nor2_1 U20711 ( .A(n24009), .B(n23972), .Y(n13940) );
  nor2_1 U20712 ( .A(n10626), .B(n23972), .Y(n13931) );
  nor2_1 U20713 ( .A(n1678), .B(n24008), .Y(n13939) );
  o21ai_0 U20714 ( .A1(n20559), .A2(n16838), .B1(n16840), .Y(n20401) );
  xor2_1 U20715 ( .A(n16829), .B(n20560), .X(n16840) );
  nor2_1 U20716 ( .A(n18256), .B(n10609), .Y(n20560) );
  a21oi_1 U20717 ( .A1(n16835), .A2(n16833), .B1(n20561), .Y(n16838) );
  inv_1 U20718 ( .A(n16834), .Y(n20561) );
  xor2_1 U20719 ( .A(n19375), .B(n20562), .X(n16834) );
  nor2_1 U20720 ( .A(n15880), .B(n18439), .Y(n20562) );
  inv_1 U20721 ( .A(n17550), .Y(n19375) );
  nand2_1 U20722 ( .A(n20563), .B(n16826), .Y(n16833) );
  inv_1 U20723 ( .A(n16836), .Y(n16826) );
  xor2_1 U20724 ( .A(n18680), .B(n20564), .X(n16836) );
  and2_0 U20725 ( .A(n18446), .B(n12331), .X(n20564) );
  inv_1 U20726 ( .A(n19327), .Y(n18680) );
  xor2_1 U20727 ( .A(n16825), .B(n19327), .X(n20563) );
  nor3_1 U20728 ( .A(n19683), .B(n20447), .C(n20565), .Y(n19327) );
  inv_1 U20729 ( .A(n12385), .Y(n20447) );
  nand2_1 U20730 ( .A(n24035), .B(n12403), .Y(n12385) );
  inv_1 U20731 ( .A(n24023), .Y(n12403) );
  inv_1 U20732 ( .A(n12404), .Y(n19683) );
  nor3_1 U20733 ( .A(n16837), .B(n24019), .C(n18449), .Y(n16825) );
  xor2_1 U20734 ( .A(n20566), .B(n20567), .X(n18449) );
  xor2_1 U20735 ( .A(n20568), .B(n18840), .X(n20567) );
  nand2_1 U20736 ( .A(n13402), .B(n20569), .Y(n18840) );
  nand3_1 U20737 ( .A(n24003), .B(n13409), .C(n24020), .Y(n20569) );
  nand3_1 U20738 ( .A(n13383), .B(n13384), .C(n13387), .Y(n13402) );
  inv_1 U20739 ( .A(n19560), .Y(n13387) );
  xor2_1 U20740 ( .A(n10609), .B(n12331), .X(n20566) );
  nor2_1 U20741 ( .A(n18446), .B(n12331), .Y(n16837) );
  xnor2_1 U20742 ( .A(n20570), .B(n20571), .Y(n18446) );
  nand2_1 U20743 ( .A(n18439), .B(n15880), .Y(n16835) );
  xor2_1 U20744 ( .A(n20572), .B(n20573), .X(n18439) );
  xor2_1 U20745 ( .A(n10609), .B(n24022), .X(n20572) );
  inv_1 U20746 ( .A(n16841), .Y(n20559) );
  nand2_1 U20747 ( .A(n18256), .B(n10609), .Y(n16841) );
  xor2_1 U20748 ( .A(n20574), .B(n20575), .X(n18256) );
  xor2_1 U20749 ( .A(n24011), .B(n12333), .X(n20575) );
  xor2_1 U20750 ( .A(n20576), .B(n11570), .X(n20574) );
  a211oi_1 U20751 ( .A1(n19087), .A2(n20130), .B1(n20577), .C1(n20578), .Y(
        n11570) );
  o21ai_0 U20752 ( .A1(n16190), .A2(n10605), .B1(n16184), .Y(n20578) );
  inv_1 U20753 ( .A(n16187), .Y(n20130) );
  xor2_1 U20754 ( .A(n20579), .B(n20580), .X(n18432) );
  xor2_1 U20755 ( .A(n24011), .B(n12401), .X(n20580) );
  xor2_1 U20756 ( .A(n20581), .B(n11520), .X(n20579) );
  inv_1 U20757 ( .A(n12297), .Y(n11520) );
  inv_1 U20758 ( .A(n18426), .Y(n20403) );
  xor2_1 U20759 ( .A(n20582), .B(n20583), .X(n18426) );
  xor2_1 U20760 ( .A(n23993), .B(n12305), .X(n20583) );
  xor2_1 U20761 ( .A(n20584), .B(n18535), .X(n20582) );
  inv_1 U20762 ( .A(n11621), .Y(n18535) );
  nand2_1 U20763 ( .A(n14701), .B(n14693), .Y(n11621) );
  nand2_1 U20764 ( .A(n24040), .B(n20585), .Y(n14701) );
  xor2_1 U20765 ( .A(n20586), .B(n15988), .X(n18292) );
  xor2_1 U20766 ( .A(n12401), .B(n12388), .X(n15988) );
  inv_1 U20767 ( .A(n18420), .Y(n18241) );
  xor2_1 U20768 ( .A(n20587), .B(n20588), .X(n18420) );
  xor2_1 U20769 ( .A(n23985), .B(n12305), .X(n20588) );
  xor2_1 U20770 ( .A(n20589), .B(n20590), .X(n18296) );
  xor2_1 U20771 ( .A(n20591), .B(n16931), .X(n20589) );
  xor2_1 U20772 ( .A(n20592), .B(n20593), .X(n20420) );
  xor2_1 U20773 ( .A(n12392), .B(n19837), .X(n20593) );
  a21oi_1 U20774 ( .A1(n14693), .A2(n24040), .B1(n14661), .Y(n19837) );
  nor2_1 U20775 ( .A(n23986), .B(n24040), .Y(n14661) );
  inv_1 U20776 ( .A(n24042), .Y(n14693) );
  nand2_1 U20777 ( .A(n20594), .B(n20595), .Y(n20592) );
  inv_1 U20778 ( .A(n18223), .Y(n18222) );
  o22ai_1 U20779 ( .A1(n20596), .A2(n20597), .B1(n23981), .B2(n20598), .Y(
        n18223) );
  and2_0 U20780 ( .A(n20599), .B(n20600), .X(n20598) );
  inv_1 U20781 ( .A(n18303), .Y(n18400) );
  xor2_1 U20782 ( .A(n20601), .B(n20602), .X(n18303) );
  xor2_1 U20783 ( .A(n10606), .B(n12392), .X(n20601) );
  and2_0 U20784 ( .A(n18309), .B(n15990), .X(n20426) );
  inv_1 U20785 ( .A(n11574), .Y(n16750) );
  nand2_1 U20786 ( .A(n13401), .B(n13368), .Y(n11574) );
  nand2_1 U20787 ( .A(n23995), .B(n23979), .Y(n13368) );
  nand2_1 U20788 ( .A(n12821), .B(n13410), .Y(n13401) );
  inv_1 U20789 ( .A(n23995), .Y(n13410) );
  xnor2_1 U20790 ( .A(n20603), .B(n15910), .Y(n18309) );
  xor2_1 U20791 ( .A(n12340), .B(n12393), .X(n15910) );
  inv_1 U20792 ( .A(n18311), .Y(n18394) );
  xor2_1 U20793 ( .A(n20604), .B(n20605), .X(n18311) );
  inv_1 U20794 ( .A(n24045), .Y(n14685) );
  inv_1 U20795 ( .A(n18383), .Y(n18320) );
  xor2_1 U20796 ( .A(n20606), .B(n20607), .X(n18383) );
  xor2_1 U20797 ( .A(n23958), .B(n12319), .X(n20607) );
  xor2_1 U20798 ( .A(n20608), .B(n20609), .X(n18371) );
  xor2_1 U20799 ( .A(n23948), .B(n12319), .X(n20609) );
  inv_1 U20800 ( .A(n17620), .Y(n18118) );
  o221ai_1 U20801 ( .A1(n10615), .A2(n16175), .B1(n10605), .B2(n19911), .C1(
        n16184), .Y(n17620) );
  inv_1 U20802 ( .A(n18377), .Y(n18373) );
  xor2_1 U20803 ( .A(n20610), .B(n20611), .X(n18377) );
  xor2_1 U20804 ( .A(n23953), .B(n12302), .X(n20611) );
  xor2_1 U20805 ( .A(n20612), .B(n11710), .X(n20610) );
  nor2_1 U20806 ( .A(n20613), .B(n19238), .Y(n11710) );
  nor2_1 U20807 ( .A(n13957), .B(n23992), .Y(n19238) );
  inv_1 U20808 ( .A(n19855), .Y(n13957) );
  nor2_1 U20809 ( .A(n19236), .B(n23990), .Y(n19855) );
  mux2_1 U20810 ( .A0(n13938), .A1(n13952), .S(n23990), .X(n20613) );
  nor2_1 U20811 ( .A(n18368), .B(n12302), .Y(n20444) );
  inv_1 U20812 ( .A(n18336), .Y(n18368) );
  xor2_1 U20813 ( .A(n20614), .B(n20615), .X(n18336) );
  xor2_1 U20814 ( .A(n23948), .B(n12299), .X(n20615) );
  xor2_1 U20815 ( .A(n20616), .B(n11650), .X(n20614) );
  nand3_1 U20816 ( .A(n19744), .B(n16147), .C(n20617), .Y(n11292) );
  a22oi_1 U20817 ( .A1(n19747), .A2(n19235), .B1(n13886), .B2(n13928), .Y(
        n20617) );
  inv_1 U20818 ( .A(n13930), .Y(n13886) );
  nand2_1 U20819 ( .A(n23970), .B(n23990), .Y(n13930) );
  inv_1 U20820 ( .A(n13950), .Y(n19747) );
  nand2_1 U20821 ( .A(n23990), .B(n19236), .Y(n13950) );
  inv_1 U20822 ( .A(n23970), .Y(n19236) );
  nand2_1 U20823 ( .A(n13821), .B(n13924), .Y(n16147) );
  nor2_1 U20824 ( .A(n23990), .B(n23970), .Y(n13924) );
  nand2_1 U20825 ( .A(n13938), .B(n23970), .Y(n19744) );
  inv_1 U20826 ( .A(n19234), .Y(n13938) );
  nand2_1 U20827 ( .A(n23991), .B(n13928), .Y(n19234) );
  xnor2_1 U20828 ( .A(n20618), .B(n15947), .Y(n18193) );
  xor2_1 U20829 ( .A(n20619), .B(n20620), .X(n18345) );
  xor2_1 U20830 ( .A(n12320), .B(n12299), .X(n20620) );
  xor2_1 U20831 ( .A(n20621), .B(n20622), .X(n18346) );
  xor2_1 U20832 ( .A(n23938), .B(n18477), .X(n20622) );
  nand2_1 U20833 ( .A(n20623), .B(n20624), .Y(n20621) );
  xnor2_1 U20834 ( .A(n20625), .B(n20626), .Y(n18178) );
  xor2_1 U20835 ( .A(n20627), .B(n19241), .X(n20626) );
  inv_1 U20836 ( .A(n12817), .Y(n19241) );
  o21ai_0 U20837 ( .A1(n12223), .A2(n20258), .B1(n20628), .Y(n12817) );
  xor2_1 U20838 ( .A(n20629), .B(n20630), .X(n18350) );
  xor2_1 U20839 ( .A(n23949), .B(n23938), .X(n20630) );
  xor2_1 U20840 ( .A(n16934), .B(n20631), .X(n20629) );
  nand3_1 U20841 ( .A(n12409), .B(n12404), .C(n12424), .Y(n16934) );
  nand2_1 U20842 ( .A(n12422), .B(n24035), .Y(n12424) );
  nor2_1 U20843 ( .A(n20258), .B(n24023), .Y(n12422) );
  nand2_1 U20844 ( .A(n12223), .B(n20258), .Y(n12404) );
  nand2_1 U20845 ( .A(n20565), .B(n12410), .Y(n12409) );
  nor2_1 U20846 ( .A(n20258), .B(n12383), .Y(n20565) );
  inv_1 U20847 ( .A(n24031), .Y(n20258) );
  xnor2_1 U20848 ( .A(n20632), .B(n16007), .Y(n18163) );
  xor2_1 U20849 ( .A(n20633), .B(n12984), .X(n20632) );
  inv_1 U20850 ( .A(n12726), .Y(n12984) );
  nand2_1 U20851 ( .A(n20634), .B(n19911), .Y(n12726) );
  o21ai_0 U20852 ( .A1(n24004), .A2(n20543), .B1(n19814), .Y(n20634) );
  nand2_1 U20853 ( .A(n24004), .B(n16187), .Y(n19814) );
  nand2_1 U20854 ( .A(n24006), .B(n24007), .Y(n16187) );
  inv_1 U20855 ( .A(n16190), .Y(n20543) );
  nand2_1 U20856 ( .A(n20628), .B(n20186), .Y(n17550) );
  nand2_1 U20857 ( .A(n12222), .B(n12410), .Y(n20186) );
  inv_1 U20858 ( .A(n12334), .Y(n12222) );
  nand2_1 U20859 ( .A(n24023), .B(n24031), .Y(n12334) );
  a21oi_1 U20860 ( .A1(n12223), .A2(n24023), .B1(n19684), .Y(n20628) );
  nor3_1 U20861 ( .A(n24025), .B(n24031), .C(n24023), .Y(n19684) );
  inv_1 U20862 ( .A(n12335), .Y(n12223) );
  nand2_1 U20863 ( .A(n12383), .B(n12410), .Y(n12335) );
  inv_1 U20864 ( .A(n24035), .Y(n12410) );
  inv_1 U20865 ( .A(n24025), .Y(n12383) );
  inv_1 U20866 ( .A(n18157), .Y(n20307) );
  xnor2_1 U20867 ( .A(n20188), .B(n20635), .Y(n18157) );
  mux2i_1 U20868 ( .A0(n20636), .A1(n20637), .S(n18397), .Y(n20635) );
  inv_1 U20869 ( .A(n17611), .Y(n18397) );
  nand3_1 U20870 ( .A(n20638), .B(n16188), .C(n20639), .Y(n17611) );
  a22oi_1 U20871 ( .A1(n18843), .A2(n20640), .B1(n20360), .B2(n16134), .Y(
        n20639) );
  o21ai_0 U20872 ( .A1(n23976), .A2(n23974), .B1(n16164), .Y(n20640) );
  nand2_1 U20873 ( .A(n23976), .B(n23974), .Y(n16164) );
  inv_1 U20874 ( .A(n20358), .Y(n18843) );
  nand2_1 U20875 ( .A(n16124), .B(n23975), .Y(n20358) );
  inv_1 U20876 ( .A(n16176), .Y(n16124) );
  nand2_1 U20877 ( .A(n23977), .B(n23978), .Y(n16176) );
  nand2_1 U20878 ( .A(n20360), .B(n16163), .Y(n16188) );
  inv_1 U20879 ( .A(n23975), .Y(n16163) );
  inv_1 U20880 ( .A(n20092), .Y(n20360) );
  nand2_1 U20881 ( .A(n23976), .B(n19414), .Y(n20092) );
  inv_1 U20882 ( .A(n23974), .Y(n19414) );
  o21ai_0 U20883 ( .A1(n16134), .A2(n16071), .B1(n20462), .Y(n20638) );
  inv_1 U20884 ( .A(n16178), .Y(n20462) );
  nand2_1 U20885 ( .A(n19955), .B(n23975), .Y(n16178) );
  inv_1 U20886 ( .A(n18845), .Y(n19955) );
  nand2_1 U20887 ( .A(n23974), .B(n19415), .Y(n18845) );
  inv_1 U20888 ( .A(n23976), .Y(n19415) );
  inv_1 U20889 ( .A(n16158), .Y(n16071) );
  nand2_1 U20890 ( .A(n23977), .B(n19407), .Y(n16158) );
  nor2_1 U20891 ( .A(n19407), .B(n23977), .Y(n16134) );
  inv_1 U20892 ( .A(n23978), .Y(n19407) );
  o22ai_1 U20893 ( .A1(n20641), .A2(n10826), .B1(n20642), .B2(n10607), .Y(
        n20637) );
  nor2_1 U20894 ( .A(n12380), .B(n20633), .Y(n20642) );
  inv_1 U20895 ( .A(n12380), .Y(n10826) );
  and2_0 U20896 ( .A(n16007), .B(n20641), .X(n20636) );
  inv_1 U20897 ( .A(n20633), .Y(n20641) );
  o22ai_1 U20898 ( .A1(n23938), .A2(n20631), .B1(n20643), .B2(n16015), .Y(
        n20633) );
  inv_1 U20899 ( .A(n23949), .Y(n16015) );
  and2_0 U20900 ( .A(n20631), .B(n23938), .X(n20643) );
  xnor2_1 U20901 ( .A(n20644), .B(n23979), .Y(n20631) );
  mux2i_1 U20902 ( .A0(n20645), .A1(n20646), .S(n10958), .Y(n20644) );
  inv_1 U20903 ( .A(n16904), .Y(n10958) );
  a21oi_1 U20904 ( .A1(n20647), .A2(n15953), .B1(n20648), .Y(n20646) );
  a21oi_1 U20905 ( .A1(n20627), .A2(n12320), .B1(n23950), .Y(n20648) );
  nand2_1 U20906 ( .A(n20627), .B(n20625), .Y(n20645) );
  xor2_1 U20907 ( .A(n10607), .B(n15953), .X(n20625) );
  inv_1 U20908 ( .A(n20647), .Y(n20627) );
  o21ai_0 U20909 ( .A1(n20649), .A2(n16013), .B1(n20624), .Y(n20647) );
  o221ai_1 U20910 ( .A1(n12320), .A2(n20650), .B1(n12299), .B2(n20619), .C1(
        n23951), .Y(n20624) );
  nor2_1 U20911 ( .A(n15955), .B(n20651), .Y(n20650) );
  inv_1 U20912 ( .A(n23938), .Y(n16013) );
  inv_1 U20913 ( .A(n20623), .Y(n20649) );
  o221ai_1 U20914 ( .A1(n20652), .A2(n15953), .B1(n15955), .B2(n20651), .C1(
        n20209), .Y(n20623) );
  inv_1 U20915 ( .A(n20619), .Y(n20651) );
  inv_1 U20916 ( .A(n12320), .Y(n15953) );
  nor2_1 U20917 ( .A(n12299), .B(n20619), .Y(n20652) );
  mux2i_1 U20918 ( .A0(n20653), .A1(n20654), .S(n24045), .Y(n20619) );
  o22ai_1 U20919 ( .A1(n20618), .A2(n16611), .B1(n20655), .B2(n20209), .Y(
        n20654) );
  nor2_1 U20920 ( .A(n23953), .B(n20656), .Y(n20655) );
  inv_1 U20921 ( .A(n23953), .Y(n16611) );
  nand2_1 U20922 ( .A(n20656), .B(n15947), .Y(n20653) );
  o21ai_0 U20923 ( .A1(n23953), .A2(n20209), .B1(n15956), .Y(n15947) );
  nand2_1 U20924 ( .A(n23953), .B(n20209), .Y(n15956) );
  inv_1 U20925 ( .A(n23951), .Y(n20209) );
  inv_1 U20926 ( .A(n20618), .Y(n20656) );
  xor2_1 U20927 ( .A(n20657), .B(n18077), .X(n20618) );
  inv_1 U20928 ( .A(n10879), .Y(n18077) );
  o211ai_1 U20929 ( .A1(n23962), .A2(n20658), .B1(n20659), .C1(n20660), .Y(
        n10879) );
  mux2i_1 U20930 ( .A0(n16087), .A1(n16100), .S(n23961), .Y(n20660) );
  inv_1 U20931 ( .A(n16140), .Y(n16100) );
  nand2_1 U20932 ( .A(n23963), .B(n20480), .Y(n16140) );
  inv_1 U20933 ( .A(n23960), .Y(n20480) );
  inv_1 U20934 ( .A(n20052), .Y(n16087) );
  nand2_1 U20935 ( .A(n23960), .B(n20281), .Y(n20052) );
  inv_1 U20936 ( .A(n23963), .Y(n20281) );
  mux2i_1 U20937 ( .A0(n20661), .A1(n16137), .S(n23960), .Y(n20659) );
  and2_0 U20938 ( .A(n16101), .B(n23962), .X(n16137) );
  nor2_1 U20939 ( .A(n10616), .B(n23961), .Y(n16101) );
  nor2_1 U20940 ( .A(n16155), .B(n16189), .Y(n20661) );
  nand2_1 U20941 ( .A(n23964), .B(n23961), .Y(n16189) );
  inv_1 U20942 ( .A(n23962), .Y(n16155) );
  mux2i_1 U20943 ( .A0(n10616), .A1(n23961), .S(n23963), .Y(n20658) );
  o22ai_1 U20944 ( .A1(n20662), .A2(n15955), .B1(n23948), .B2(n20663), .Y(
        n20657) );
  nor2_1 U20945 ( .A(n12299), .B(n20616), .Y(n20663) );
  inv_1 U20946 ( .A(n12299), .Y(n15955) );
  inv_1 U20947 ( .A(n20616), .Y(n20662) );
  o22ai_1 U20948 ( .A1(n15931), .A2(n20612), .B1(n23953), .B2(n20664), .Y(
        n20616) );
  and2_0 U20949 ( .A(n20612), .B(n15931), .X(n20664) );
  o22ai_1 U20950 ( .A1(n12319), .A2(n20608), .B1(n23948), .B2(n20665), .Y(
        n20612) );
  nor2_1 U20951 ( .A(n16524), .B(n20666), .Y(n20665) );
  inv_1 U20952 ( .A(n20608), .Y(n20666) );
  xor2_1 U20953 ( .A(n11489), .B(n20667), .X(n20608) );
  mux2i_1 U20954 ( .A0(n20668), .A1(n20669), .S(n18477), .Y(n20667) );
  o22ai_1 U20955 ( .A1(n20507), .A2(n15931), .B1(n23959), .B2(n20670), .Y(
        n20669) );
  nor2_1 U20956 ( .A(n12302), .B(n20671), .Y(n20670) );
  nor2_1 U20957 ( .A(n20508), .B(n20671), .Y(n20668) );
  inv_1 U20958 ( .A(n20507), .Y(n20671) );
  xor2_1 U20959 ( .A(n20672), .B(n17036), .X(n20507) );
  inv_1 U20960 ( .A(n18213), .Y(n17036) );
  nand2_1 U20961 ( .A(n20673), .B(n20674), .Y(n18213) );
  mux2i_1 U20962 ( .A0(n13397), .A1(n24020), .S(n13400), .Y(n20673) );
  inv_1 U20963 ( .A(n13367), .Y(n13400) );
  nand2_1 U20964 ( .A(n24002), .B(n19562), .Y(n13367) );
  nor2_1 U20965 ( .A(n13383), .B(n24020), .Y(n13397) );
  o22ai_1 U20966 ( .A1(n16524), .A2(n20675), .B1(n20676), .B2(n18413), .Y(
        n20672) );
  nor2_1 U20967 ( .A(n12319), .B(n20606), .Y(n20676) );
  inv_1 U20968 ( .A(n20606), .Y(n20675) );
  xor2_1 U20969 ( .A(n20677), .B(n18477), .X(n20606) );
  inv_1 U20970 ( .A(n17174), .Y(n18477) );
  o22ai_1 U20971 ( .A1(n13336), .A2(n13408), .B1(n13382), .B2(n13403), .Y(
        n17174) );
  nand2_1 U20972 ( .A(n10622), .B(n13398), .Y(n13403) );
  o22ai_1 U20973 ( .A1(n12393), .A2(n20513), .B1(n23959), .B2(n20678), .Y(
        n20677) );
  and2_0 U20974 ( .A(n12393), .B(n20513), .X(n20678) );
  mux2i_1 U20975 ( .A0(n20679), .A1(n20680), .S(n18068), .Y(n20513) );
  inv_1 U20976 ( .A(n19338), .Y(n18068) );
  o21ai_0 U20977 ( .A1(n19087), .A2(n16190), .B1(n20681), .Y(n19338) );
  mux2i_1 U20978 ( .A0(n20577), .A1(n20682), .S(n20131), .Y(n20681) );
  nor2_1 U20979 ( .A(n10605), .B(n19088), .Y(n20682) );
  nor2_1 U20980 ( .A(n19088), .B(n24004), .Y(n20577) );
  o22ai_1 U20981 ( .A1(n20604), .A2(n18413), .B1(n20683), .B2(n10606), .Y(
        n20680) );
  nor2_1 U20982 ( .A(n23958), .B(n20684), .Y(n20683) );
  nand2_1 U20983 ( .A(n20684), .B(n20605), .Y(n20679) );
  o21ai_0 U20984 ( .A1(n1965), .A2(n18413), .B1(n15909), .Y(n20605) );
  nand2_1 U20985 ( .A(n1965), .B(n18413), .Y(n15909) );
  inv_1 U20986 ( .A(n23958), .Y(n18413) );
  inv_1 U20987 ( .A(n20604), .Y(n20684) );
  xor2_1 U20988 ( .A(n20685), .B(n17765), .X(n20604) );
  a211oi_1 U20989 ( .A1(n13922), .A2(n13921), .B1(n13884), .C1(n13725), .Y(
        n17765) );
  and2_0 U20990 ( .A(n13927), .B(n13916), .X(n13725) );
  inv_1 U20991 ( .A(n13762), .Y(n13884) );
  nand2_1 U20992 ( .A(n13867), .B(n13915), .Y(n13762) );
  o22ai_1 U20993 ( .A1(n20686), .A2(n16510), .B1(n20687), .B2(n15902), .Y(
        n20685) );
  inv_1 U20994 ( .A(n12393), .Y(n15902) );
  nor2_1 U20995 ( .A(n12340), .B(n20603), .Y(n20687) );
  inv_1 U20996 ( .A(n20603), .Y(n20686) );
  o22ai_1 U20997 ( .A1(n15990), .A2(n20602), .B1(n1965), .B2(n20688), .Y(
        n20603) );
  and2_0 U20998 ( .A(n15990), .B(n20602), .X(n20688) );
  xnor2_1 U20999 ( .A(n20689), .B(n16829), .Y(n20602) );
  inv_1 U21000 ( .A(n17976), .Y(n16829) );
  o221ai_1 U21001 ( .A1(n23999), .A2(n19967), .B1(n19395), .B2(n13947), .C1(
        n19396), .Y(n17976) );
  nand2_1 U21002 ( .A(n13927), .B(n19968), .Y(n19396) );
  nor2_1 U21003 ( .A(n13921), .B(n13916), .Y(n19967) );
  nand2_1 U21004 ( .A(n20600), .B(n20597), .Y(n20689) );
  nand2_1 U21005 ( .A(n23981), .B(n20599), .Y(n20597) );
  nand2_1 U21006 ( .A(n20690), .B(n16510), .Y(n20599) );
  inv_1 U21007 ( .A(n20596), .Y(n20600) );
  nor2_1 U21008 ( .A(n16510), .B(n20690), .Y(n20596) );
  a21oi_1 U21009 ( .A1(n20594), .A2(n12392), .B1(n20691), .Y(n20690) );
  inv_1 U21010 ( .A(n20595), .Y(n20691) );
  o211ai_1 U21011 ( .A1(n15999), .A2(n20692), .B1(n20693), .C1(n15992), .Y(
        n20595) );
  o21ai_0 U21012 ( .A1(n23981), .A2(n20533), .B1(n23987), .Y(n20693) );
  o211ai_1 U21013 ( .A1(n23981), .A2(n20533), .B1(n20694), .C1(n12394), .Y(
        n20594) );
  o21ai_0 U21014 ( .A1(n15999), .A2(n20692), .B1(n16453), .Y(n20694) );
  inv_1 U21015 ( .A(n20533), .Y(n20692) );
  inv_1 U21016 ( .A(n23981), .Y(n15999) );
  xnor2_1 U21017 ( .A(n16931), .B(n20695), .Y(n20533) );
  mux2i_1 U21018 ( .A0(n20696), .A1(n20697), .S(n11650), .Y(n20695) );
  inv_1 U21019 ( .A(n17955), .Y(n11650) );
  o32ai_1 U21020 ( .A1(n20698), .A2(n20131), .A3(n16116), .B1(n24006), .B2(
        n16183), .Y(n17955) );
  inv_1 U21021 ( .A(n16141), .Y(n16116) );
  nand2_1 U21022 ( .A(n24004), .B(n19087), .Y(n16141) );
  inv_1 U21023 ( .A(n19911), .Y(n20131) );
  o21ai_0 U21024 ( .A1(n16181), .A2(n16175), .B1(n16159), .Y(n20698) );
  nand2_1 U21025 ( .A(n24005), .B(n10605), .Y(n16159) );
  inv_1 U21026 ( .A(n16174), .Y(n16181) );
  nand2_1 U21027 ( .A(n24006), .B(n10615), .Y(n16174) );
  and2_0 U21028 ( .A(n20590), .B(n20591), .X(n20697) );
  xor2_1 U21029 ( .A(n18262), .B(n15992), .X(n20590) );
  o22ai_1 U21030 ( .A1(n20591), .A2(n15992), .B1(n20699), .B2(n18262), .Y(
        n20696) );
  nor2_1 U21031 ( .A(n12394), .B(n20700), .Y(n20699) );
  inv_1 U21032 ( .A(n20591), .Y(n20700) );
  inv_1 U21033 ( .A(n12394), .Y(n15992) );
  xor2_1 U21034 ( .A(n16666), .B(n20701), .X(n20591) );
  mux2i_1 U21035 ( .A0(n20702), .A1(n20703), .S(n18999), .Y(n20701) );
  inv_1 U21036 ( .A(n12924), .Y(n18999) );
  nand4_1 U21037 ( .A(n13937), .B(n13934), .C(n13961), .D(n20704), .Y(n12924)
         );
  a22oi_1 U21038 ( .A1(n13922), .A2(n19968), .B1(n13916), .B2(n10621), .Y(
        n20704) );
  inv_1 U21039 ( .A(n13948), .Y(n13916) );
  nand2_1 U21040 ( .A(n19395), .B(n19968), .Y(n13948) );
  inv_1 U21041 ( .A(n24000), .Y(n19395) );
  inv_1 U21042 ( .A(n13947), .Y(n13922) );
  nand2_1 U21043 ( .A(n23999), .B(n10621), .Y(n13947) );
  nand2_1 U21044 ( .A(n13867), .B(n13927), .Y(n13961) );
  nor2_1 U21045 ( .A(n10621), .B(n23999), .Y(n13927) );
  inv_1 U21046 ( .A(n19970), .Y(n13867) );
  nand2_1 U21047 ( .A(n24000), .B(n19968), .Y(n19970) );
  nand2_1 U21048 ( .A(n13921), .B(n13868), .Y(n13934) );
  nor2_1 U21049 ( .A(n23998), .B(n23999), .Y(n13868) );
  inv_1 U21050 ( .A(n13960), .Y(n13921) );
  nand2_1 U21051 ( .A(n24001), .B(n24000), .Y(n13960) );
  nand2_1 U21052 ( .A(n13915), .B(n13926), .Y(n13937) );
  nor2_1 U21053 ( .A(n19968), .B(n24000), .Y(n13926) );
  inv_1 U21054 ( .A(n24001), .Y(n19968) );
  nor2_1 U21055 ( .A(n19890), .B(n10621), .Y(n13915) );
  inv_1 U21056 ( .A(n23999), .Y(n19890) );
  o22ai_1 U21057 ( .A1(n12388), .A2(n20705), .B1(n20706), .B2(n16453), .Y(
        n20703) );
  nor2_1 U21058 ( .A(n20546), .B(n15970), .Y(n20706) );
  inv_1 U21059 ( .A(n20546), .Y(n20705) );
  nor2_1 U21060 ( .A(n20546), .B(n20544), .Y(n20702) );
  xor2_1 U21061 ( .A(n16453), .B(n15970), .X(n20544) );
  inv_1 U21062 ( .A(n12388), .Y(n15970) );
  inv_1 U21063 ( .A(n23987), .Y(n16453) );
  a21oi_1 U21064 ( .A1(n20707), .A2(n12305), .B1(n20708), .Y(n20546) );
  a21oi_1 U21065 ( .A1(n15972), .A2(n20587), .B1(n18262), .Y(n20708) );
  inv_1 U21066 ( .A(n23985), .Y(n18262) );
  inv_1 U21067 ( .A(n20707), .Y(n20587) );
  o22ai_1 U21068 ( .A1(n12388), .A2(n20586), .B1(n12401), .B2(n20709), .Y(
        n20707) );
  and2_0 U21069 ( .A(n20586), .B(n12388), .X(n20709) );
  o22ai_1 U21070 ( .A1(n15972), .A2(n20584), .B1(n23993), .B2(n20710), .Y(
        n20586) );
  and2_0 U21071 ( .A(n20584), .B(n15972), .X(n20710) );
  o22ai_1 U21072 ( .A1(n18463), .A2(n20581), .B1(n20711), .B2(n10608), .Y(
        n20584) );
  and2_0 U21073 ( .A(n18463), .B(n20581), .X(n20711) );
  xor2_1 U21074 ( .A(n20712), .B(n10919), .X(n20581) );
  o221ai_1 U21075 ( .A1(n19087), .A2(n16190), .B1(n24004), .B2(n19911), .C1(
        n20713), .Y(n10919) );
  a21oi_1 U21076 ( .A1(n16093), .A2(n24006), .B1(n20714), .Y(n20713) );
  inv_1 U21077 ( .A(n16184), .Y(n20714) );
  nand2_1 U21078 ( .A(n16183), .B(n19088), .Y(n16184) );
  inv_1 U21079 ( .A(n16175), .Y(n16183) );
  nand2_1 U21080 ( .A(n24005), .B(n24004), .Y(n16175) );
  inv_1 U21081 ( .A(n16177), .Y(n16093) );
  nand2_1 U21082 ( .A(n10605), .B(n19087), .Y(n16177) );
  nand2_1 U21083 ( .A(n19087), .B(n10615), .Y(n19911) );
  nand2_1 U21084 ( .A(n19088), .B(n10615), .Y(n16190) );
  inv_1 U21085 ( .A(n24006), .Y(n19088) );
  inv_1 U21086 ( .A(n24005), .Y(n19087) );
  mux2i_1 U21087 ( .A0(n20715), .A1(n20716), .S(n12942), .Y(n20712) );
  a21oi_1 U21088 ( .A1(n13821), .A2(n23990), .B1(n13952), .Y(n12942) );
  nor3_1 U21089 ( .A(n13929), .B(n23970), .C(n13928), .Y(n13952) );
  inv_1 U21090 ( .A(n19235), .Y(n13821) );
  nand2_1 U21091 ( .A(n13929), .B(n13928), .Y(n19235) );
  inv_1 U21092 ( .A(n23992), .Y(n13928) );
  inv_1 U21093 ( .A(n23991), .Y(n13929) );
  o22ai_1 U21094 ( .A1(n20717), .A2(n15913), .B1(n23993), .B2(n20718), .Y(
        n20716) );
  nor2_1 U21095 ( .A(n24022), .B(n20558), .Y(n20718) );
  or2_0 U21096 ( .A(n20557), .B(n20717), .X(n20715) );
  inv_1 U21097 ( .A(n20558), .Y(n20717) );
  o22ai_1 U21098 ( .A1(n12333), .A2(n20719), .B1(n24011), .B2(n20720), .Y(
        n20558) );
  nor2_1 U21099 ( .A(n20576), .B(n15920), .Y(n20720) );
  inv_1 U21100 ( .A(n20576), .Y(n20719) );
  xor2_1 U21101 ( .A(n16904), .B(n20721), .X(n20576) );
  a21oi_1 U21102 ( .A1(n20573), .A2(n10609), .B1(n20722), .Y(n20721) );
  inv_1 U21103 ( .A(n20723), .Y(n20722) );
  o21ai_0 U21104 ( .A1(n10609), .A2(n20573), .B1(n24022), .Y(n20723) );
  mux2i_1 U21105 ( .A0(n20724), .A1(n20725), .S(n16843), .Y(n20573) );
  nand2_1 U21106 ( .A(n13381), .B(n20726), .Y(n16843) );
  nand3_1 U21107 ( .A(n13408), .B(n10622), .C(n13382), .Y(n20726) );
  o22ai_1 U21108 ( .A1(n15880), .A2(n20570), .B1(n20727), .B2(n15920), .Y(
        n20725) );
  inv_1 U21109 ( .A(n12333), .Y(n15920) );
  nor2_1 U21110 ( .A(n20728), .B(n12408), .Y(n20727) );
  nand2_1 U21111 ( .A(n20728), .B(n20571), .Y(n20724) );
  xor2_1 U21112 ( .A(n12408), .B(n12333), .X(n20571) );
  inv_1 U21113 ( .A(n20570), .Y(n20728) );
  o22ai_1 U21114 ( .A1(n12331), .A2(n20729), .B1(n20730), .B2(n10609), .Y(
        n20570) );
  nor2_1 U21115 ( .A(n20568), .B(n18455), .Y(n20730) );
  inv_1 U21116 ( .A(n20568), .Y(n20729) );
  o221ai_1 U21117 ( .A1(n20731), .A2(n18462), .B1(n18464), .B2(n15880), .C1(
        n20732), .Y(n20568) );
  nand2_1 U21118 ( .A(n15895), .B(n19009), .Y(n20732) );
  inv_1 U21119 ( .A(n17340), .Y(n19009) );
  o21ai_0 U21120 ( .A1(n12408), .A2(n18462), .B1(n15884), .Y(n15895) );
  nand2_1 U21121 ( .A(n12408), .B(n18462), .Y(n15884) );
  inv_1 U21122 ( .A(n12408), .Y(n15880) );
  inv_1 U21123 ( .A(n20124), .Y(n18464) );
  inv_1 U21124 ( .A(n24019), .Y(n18462) );
  a21oi_1 U21125 ( .A1(n12408), .A2(n17340), .B1(n20124), .Y(n20731) );
  xnor2_1 U21126 ( .A(n18184), .B(n16842), .Y(n20124) );
  inv_1 U21127 ( .A(n17967), .Y(n16842) );
  nand2_1 U21128 ( .A(n24019), .B(n18455), .Y(n17967) );
  inv_1 U21129 ( .A(n12331), .Y(n18455) );
  nand2_1 U21130 ( .A(n19530), .B(n12425), .Y(n18184) );
  nand2_1 U21131 ( .A(n19531), .B(n24026), .Y(n12425) );
  nor2_1 U21132 ( .A(n24032), .B(n24033), .Y(n19531) );
  inv_1 U21133 ( .A(n20733), .Y(n19530) );
  o21ai_0 U21134 ( .A1(n12423), .A2(n19529), .B1(n20336), .Y(n20733) );
  nand2_1 U21135 ( .A(n12431), .B(n12384), .Y(n20336) );
  nor2_1 U21136 ( .A(n12405), .B(n24026), .Y(n12431) );
  nand2_1 U21137 ( .A(n24033), .B(n19528), .Y(n12405) );
  inv_1 U21138 ( .A(n24032), .Y(n19528) );
  nand2_1 U21139 ( .A(n11801), .B(n12406), .Y(n19529) );
  inv_1 U21140 ( .A(n24026), .Y(n12406) );
  inv_1 U21141 ( .A(n12384), .Y(n11801) );
  nand2_1 U21142 ( .A(n24033), .B(n24032), .Y(n12423) );
  nor3_1 U21143 ( .A(n19805), .B(n20734), .C(n20735), .Y(n17340) );
  o32ai_1 U21144 ( .A1(n14687), .A2(n24047), .A3(n20252), .B1(n14696), .B2(
        n14702), .Y(n20735) );
  nand2_1 U21145 ( .A(n24038), .B(n10636), .Y(n14687) );
  mux2i_1 U21146 ( .A0(n14663), .A1(n14673), .S(n24038), .Y(n20734) );
  nand2_1 U21147 ( .A(n19671), .B(n24046), .Y(n14673) );
  inv_1 U21148 ( .A(n14696), .Y(n19671) );
  nand2_1 U21149 ( .A(n24047), .B(n20252), .Y(n14696) );
  inv_1 U21150 ( .A(n24017), .Y(n20252) );
  nand3_1 U21151 ( .A(n24046), .B(n14676), .C(n24017), .Y(n14663) );
  inv_1 U21152 ( .A(n24047), .Y(n14676) );
  o22ai_1 U21153 ( .A1(n14707), .A2(n14699), .B1(n20736), .B2(n14702), .Y(
        n19805) );
  nand2_1 U21154 ( .A(n20033), .B(n10636), .Y(n14702) );
  inv_1 U21155 ( .A(n24038), .Y(n20033) );
  a21oi_1 U21156 ( .A1(n24017), .A2(n24046), .B1(n19146), .Y(n20736) );
  nor2_1 U21157 ( .A(n24017), .B(n24046), .Y(n19146) );
  nand2_1 U21158 ( .A(n14675), .B(n24047), .Y(n14699) );
  inv_1 U21159 ( .A(n14698), .Y(n14675) );
  nand2_1 U21160 ( .A(n24017), .B(n20030), .Y(n14698) );
  inv_1 U21161 ( .A(n24046), .Y(n20030) );
  nand2_1 U21162 ( .A(n24039), .B(n24038), .Y(n14707) );
  o21ai_0 U21163 ( .A1(n19560), .A2(n13384), .B1(n20674), .Y(n16904) );
  mux2i_1 U21164 ( .A0(n13385), .A1(n24002), .S(n13386), .Y(n20674) );
  inv_1 U21165 ( .A(n13369), .Y(n13386) );
  nand2_1 U21166 ( .A(n24020), .B(n13383), .Y(n13369) );
  inv_1 U21167 ( .A(n24003), .Y(n13383) );
  nor2_1 U21168 ( .A(n19562), .B(n24002), .Y(n13385) );
  inv_1 U21169 ( .A(n24020), .Y(n13384) );
  nand2_1 U21170 ( .A(n13409), .B(n19562), .Y(n19560) );
  inv_1 U21171 ( .A(n24021), .Y(n19562) );
  inv_1 U21172 ( .A(n24002), .Y(n13409) );
  xor2_1 U21173 ( .A(n10775), .B(n15913), .X(n20557) );
  inv_1 U21174 ( .A(n24022), .Y(n15913) );
  inv_1 U21175 ( .A(n23993), .Y(n10775) );
  inv_1 U21176 ( .A(n12401), .Y(n18463) );
  inv_1 U21177 ( .A(n12305), .Y(n15972) );
  o21ai_0 U21178 ( .A1(n24042), .A2(n20585), .B1(n14705), .Y(n16666) );
  inv_1 U21179 ( .A(n14683), .Y(n14705) );
  nor2_1 U21180 ( .A(n20585), .B(n24040), .Y(n14683) );
  inv_1 U21181 ( .A(n23986), .Y(n20585) );
  and3_1 U21182 ( .A(n13395), .B(n13392), .C(n20536), .X(n16931) );
  inv_1 U21183 ( .A(n20528), .Y(n20536) );
  o22ai_1 U21184 ( .A1(n23983), .A2(n13382), .B1(n10622), .B2(n13378), .Y(
        n20528) );
  nand2_1 U21185 ( .A(n24013), .B(n20529), .Y(n13378) );
  nand2_1 U21186 ( .A(n24013), .B(n24012), .Y(n13382) );
  nand2_1 U21187 ( .A(n23982), .B(n13398), .Y(n13392) );
  inv_1 U21188 ( .A(n23983), .Y(n13398) );
  nand2_1 U21189 ( .A(n13336), .B(n20068), .Y(n13395) );
  inv_1 U21190 ( .A(n13408), .Y(n20068) );
  nand2_1 U21191 ( .A(n20529), .B(n18468), .Y(n13408) );
  inv_1 U21192 ( .A(n24013), .Y(n18468) );
  inv_1 U21193 ( .A(n24012), .Y(n20529) );
  inv_1 U21194 ( .A(n13381), .Y(n13336) );
  nand2_1 U21195 ( .A(n23983), .B(n10622), .Y(n13381) );
  inv_1 U21196 ( .A(n12340), .Y(n16510) );
  inv_1 U21197 ( .A(n12392), .Y(n15990) );
  inv_1 U21198 ( .A(n12319), .Y(n16524) );
  inv_1 U21199 ( .A(n15928), .Y(n20508) );
  o21ai_0 U21200 ( .A1(n23959), .A2(n12302), .B1(n15933), .Y(n15928) );
  nand2_1 U21201 ( .A(n23959), .B(n12302), .Y(n15933) );
  nand2_1 U21202 ( .A(n23995), .B(n12821), .Y(n11489) );
  inv_1 U21203 ( .A(n23979), .Y(n12821) );
  inv_1 U21204 ( .A(n12302), .Y(n15931) );
  o21ai_0 U21205 ( .A1(n12380), .A2(n10607), .B1(n19981), .Y(n16007) );
  nand2_1 U21206 ( .A(n12380), .B(n10607), .Y(n19981) );
  nor2_1 U21207 ( .A(n20737), .B(n18765), .Y(n20188) );
  nor2_1 U21208 ( .A(n12380), .B(n23949), .Y(n18765) );
  inv_1 U21209 ( .A(n18764), .Y(n20737) );
  nand2_1 U21210 ( .A(n23949), .B(n12380), .Y(n18764) );
  o21ai_0 U21211 ( .A1(n20738), .A2(n15875), .B1(n11482), .Y(n11480) );
  or2_0 U21212 ( .A(n11402), .B(n20738), .X(n11482) );
  nand2_1 U21213 ( .A(n16951), .B(n11400), .Y(n11402) );
  nand2_1 U21214 ( .A(n15815), .B(n15718), .Y(n11400) );
  inv_1 U21215 ( .A(n11211), .Y(n15815) );
  nand2_1 U21216 ( .A(n20739), .B(n15875), .Y(n11211) );
  a21oi_1 U21217 ( .A1(n24051), .A2(n15851), .B1(n15872), .Y(n16951) );
  nor2_1 U21218 ( .A(n16206), .B(n15875), .Y(n15872) );
  nand2_1 U21219 ( .A(n24051), .B(n20739), .Y(n16206) );
  inv_1 U21220 ( .A(n24048), .Y(n20739) );
  inv_1 U21221 ( .A(n15858), .Y(n15851) );
  nand2_1 U21222 ( .A(n24048), .B(n15875), .Y(n15858) );
  inv_1 U21223 ( .A(n24054), .Y(n15875) );
  inv_1 U21224 ( .A(n11150), .Y(n20738) );
  nand2_1 U21225 ( .A(n15870), .B(n15718), .Y(n11150) );
  inv_1 U21226 ( .A(n24051), .Y(n15718) );
  inv_1 U21227 ( .A(n15859), .Y(n15870) );
  nand2_1 U21228 ( .A(n24048), .B(n24054), .Y(n15859) );
  nor2_1 U21229 ( .A(n19445), .B(n19964), .Y(n19449) );
  inv_1 U21230 ( .A(n19446), .Y(n19964) );
  nand2_1 U21231 ( .A(n12308), .B(outData[0]), .Y(n19446) );
  nor2_1 U21232 ( .A(outData[0]), .B(n12308), .Y(n19445) );
  inv_1 U21233 ( .A(n12464), .Y(outData[0]) );
endmodule

